module Sig_op6_0(
  input        clock,
  input        reset,
  input  [5:0] io_A,
  input  [5:0] io_B,
  output       io_greaterSign,
  output       io_smallerSign,
  output [3:0] io_greaterExp,
  output [4:0] io_greaterSig,
  output [7:0] io_smallerSig,
  output       io_AisNar,
  output       io_BisNar,
  output       io_AisZero,
  output       io_BisZero
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [3:0] _T_4; // @[convert.scala 19:24]
  wire [3:0] _T_5; // @[convert.scala 19:43]
  wire [3:0] _T_6; // @[convert.scala 19:39]
  wire [1:0] _T_7; // @[LZD.scala 43:32]
  wire  _T_8; // @[LZD.scala 39:14]
  wire  _T_9; // @[LZD.scala 39:21]
  wire  _T_10; // @[LZD.scala 39:30]
  wire  _T_11; // @[LZD.scala 39:27]
  wire  _T_12; // @[LZD.scala 39:25]
  wire [1:0] _T_13; // @[Cat.scala 29:58]
  wire [1:0] _T_14; // @[LZD.scala 44:32]
  wire  _T_15; // @[LZD.scala 39:14]
  wire  _T_16; // @[LZD.scala 39:21]
  wire  _T_17; // @[LZD.scala 39:30]
  wire  _T_18; // @[LZD.scala 39:27]
  wire  _T_19; // @[LZD.scala 39:25]
  wire [1:0] _T_20; // @[Cat.scala 29:58]
  wire  _T_21; // @[Shift.scala 12:21]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[LZD.scala 49:16]
  wire  _T_24; // @[LZD.scala 49:27]
  wire  _T_25; // @[LZD.scala 49:25]
  wire  _T_26; // @[LZD.scala 49:47]
  wire  _T_27; // @[LZD.scala 49:59]
  wire  _T_28; // @[LZD.scala 49:35]
  wire [2:0] _T_30; // @[Cat.scala 29:58]
  wire [2:0] _T_31; // @[convert.scala 21:22]
  wire [2:0] _T_32; // @[convert.scala 22:36]
  wire  _T_33; // @[Shift.scala 16:24]
  wire [1:0] _T_34; // @[Shift.scala 17:37]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[Shift.scala 64:52]
  wire [2:0] _T_38; // @[Cat.scala 29:58]
  wire [2:0] _T_39; // @[Shift.scala 64:27]
  wire  _T_40; // @[Shift.scala 66:70]
  wire [1:0] _T_42; // @[Shift.scala 64:52]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire [2:0] _T_44; // @[Shift.scala 64:27]
  wire [2:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_48; // @[convert.scala 25:26]
  wire [2:0] _T_50; // @[convert.scala 25:42]
  wire [3:0] _T_51; // @[Cat.scala 29:58]
  wire [4:0] _T_53; // @[convert.scala 29:56]
  wire  _T_54; // @[convert.scala 29:60]
  wire  _T_55; // @[convert.scala 29:41]
  wire  _T_58; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [3:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_67; // @[convert.scala 18:24]
  wire  _T_68; // @[convert.scala 18:40]
  wire  _T_69; // @[convert.scala 18:36]
  wire [3:0] _T_70; // @[convert.scala 19:24]
  wire [3:0] _T_71; // @[convert.scala 19:43]
  wire [3:0] _T_72; // @[convert.scala 19:39]
  wire [1:0] _T_73; // @[LZD.scala 43:32]
  wire  _T_74; // @[LZD.scala 39:14]
  wire  _T_75; // @[LZD.scala 39:21]
  wire  _T_76; // @[LZD.scala 39:30]
  wire  _T_77; // @[LZD.scala 39:27]
  wire  _T_78; // @[LZD.scala 39:25]
  wire [1:0] _T_79; // @[Cat.scala 29:58]
  wire [1:0] _T_80; // @[LZD.scala 44:32]
  wire  _T_81; // @[LZD.scala 39:14]
  wire  _T_82; // @[LZD.scala 39:21]
  wire  _T_83; // @[LZD.scala 39:30]
  wire  _T_84; // @[LZD.scala 39:27]
  wire  _T_85; // @[LZD.scala 39:25]
  wire [1:0] _T_86; // @[Cat.scala 29:58]
  wire  _T_87; // @[Shift.scala 12:21]
  wire  _T_88; // @[Shift.scala 12:21]
  wire  _T_89; // @[LZD.scala 49:16]
  wire  _T_90; // @[LZD.scala 49:27]
  wire  _T_91; // @[LZD.scala 49:25]
  wire  _T_92; // @[LZD.scala 49:47]
  wire  _T_93; // @[LZD.scala 49:59]
  wire  _T_94; // @[LZD.scala 49:35]
  wire [2:0] _T_96; // @[Cat.scala 29:58]
  wire [2:0] _T_97; // @[convert.scala 21:22]
  wire [2:0] _T_98; // @[convert.scala 22:36]
  wire  _T_99; // @[Shift.scala 16:24]
  wire [1:0] _T_100; // @[Shift.scala 17:37]
  wire  _T_101; // @[Shift.scala 12:21]
  wire  _T_102; // @[Shift.scala 64:52]
  wire [2:0] _T_104; // @[Cat.scala 29:58]
  wire [2:0] _T_105; // @[Shift.scala 64:27]
  wire  _T_106; // @[Shift.scala 66:70]
  wire [1:0] _T_108; // @[Shift.scala 64:52]
  wire [2:0] _T_109; // @[Cat.scala 29:58]
  wire [2:0] _T_110; // @[Shift.scala 64:27]
  wire [2:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_114; // @[convert.scala 25:26]
  wire [2:0] _T_116; // @[convert.scala 25:42]
  wire [3:0] _T_117; // @[Cat.scala 29:58]
  wire [4:0] _T_119; // @[convert.scala 29:56]
  wire  _T_120; // @[convert.scala 29:60]
  wire  _T_121; // @[convert.scala 29:41]
  wire  _T_124; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [3:0] decB_scale; // @[convert.scala 32:24]
  wire  aGTb; // @[Sig_op.scala 38:32]
  wire [3:0] smallerExp; // @[Sig_op.scala 42:24]
  wire [2:0] greaterFrac; // @[Sig_op.scala 43:24]
  wire [2:0] smallerFrac; // @[Sig_op.scala 44:24]
  wire  smallerZero; // @[Sig_op.scala 45:24]
  wire [3:0] _T_136; // @[Sig_op.scala 46:35]
  wire [3:0] scale_diff; // @[Sig_op.scala 46:35]
  wire  _T_137; // @[Sig_op.scala 51:53]
  wire  _T_138; // @[Sig_op.scala 51:36]
  wire [7:0] _T_141; // @[Cat.scala 29:58]
  wire [3:0] _T_142; // @[Sig_op.scala 51:124]
  wire  _T_143; // @[Shift.scala 39:24]
  wire [2:0] _T_144; // @[Shift.scala 40:44]
  wire [3:0] _T_145; // @[Shift.scala 90:30]
  wire [3:0] _T_146; // @[Shift.scala 90:48]
  wire  _T_147; // @[Shift.scala 90:57]
  wire [3:0] _GEN_0; // @[Shift.scala 90:39]
  wire [3:0] _T_148; // @[Shift.scala 90:39]
  wire  _T_149; // @[Shift.scala 12:21]
  wire  _T_150; // @[Shift.scala 12:21]
  wire [3:0] _T_152; // @[Bitwise.scala 71:12]
  wire [7:0] _T_153; // @[Cat.scala 29:58]
  wire [7:0] _T_154; // @[Shift.scala 91:22]
  wire [1:0] _T_155; // @[Shift.scala 92:77]
  wire [5:0] _T_156; // @[Shift.scala 90:30]
  wire [1:0] _T_157; // @[Shift.scala 90:48]
  wire  _T_158; // @[Shift.scala 90:57]
  wire [5:0] _GEN_1; // @[Shift.scala 90:39]
  wire [5:0] _T_159; // @[Shift.scala 90:39]
  wire  _T_160; // @[Shift.scala 12:21]
  wire  _T_161; // @[Shift.scala 12:21]
  wire [1:0] _T_163; // @[Bitwise.scala 71:12]
  wire [7:0] _T_164; // @[Cat.scala 29:58]
  wire [7:0] _T_165; // @[Shift.scala 91:22]
  wire  _T_166; // @[Shift.scala 92:77]
  wire [6:0] _T_167; // @[Shift.scala 90:30]
  wire  _T_168; // @[Shift.scala 90:48]
  wire [6:0] _GEN_2; // @[Shift.scala 90:39]
  wire [6:0] _T_170; // @[Shift.scala 90:39]
  wire  _T_172; // @[Shift.scala 12:21]
  wire [7:0] _T_173; // @[Cat.scala 29:58]
  wire [7:0] _T_174; // @[Shift.scala 91:22]
  wire [7:0] _T_177; // @[Bitwise.scala 71:12]
  wire  _T_178; // @[Sig_op.scala 57:40]
  wire [1:0] _T_179; // @[Cat.scala 29:58]
  assign _T_1 = io_A[5]; // @[convert.scala 18:24]
  assign _T_2 = io_A[4]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[4:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[3:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[3:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7 != 2'h0; // @[LZD.scala 39:14]
  assign _T_9 = _T_7[1]; // @[LZD.scala 39:21]
  assign _T_10 = _T_7[0]; // @[LZD.scala 39:30]
  assign _T_11 = ~ _T_10; // @[LZD.scala 39:27]
  assign _T_12 = _T_9 | _T_11; // @[LZD.scala 39:25]
  assign _T_13 = {_T_8,_T_12}; // @[Cat.scala 29:58]
  assign _T_14 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_15 = _T_14 != 2'h0; // @[LZD.scala 39:14]
  assign _T_16 = _T_14[1]; // @[LZD.scala 39:21]
  assign _T_17 = _T_14[0]; // @[LZD.scala 39:30]
  assign _T_18 = ~ _T_17; // @[LZD.scala 39:27]
  assign _T_19 = _T_16 | _T_18; // @[LZD.scala 39:25]
  assign _T_20 = {_T_15,_T_19}; // @[Cat.scala 29:58]
  assign _T_21 = _T_13[1]; // @[Shift.scala 12:21]
  assign _T_22 = _T_20[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21 | _T_22; // @[LZD.scala 49:16]
  assign _T_24 = ~ _T_22; // @[LZD.scala 49:27]
  assign _T_25 = _T_21 | _T_24; // @[LZD.scala 49:25]
  assign _T_26 = _T_13[0:0]; // @[LZD.scala 49:47]
  assign _T_27 = _T_20[0:0]; // @[LZD.scala 49:59]
  assign _T_28 = _T_21 ? _T_26 : _T_27; // @[LZD.scala 49:35]
  assign _T_30 = {_T_23,_T_25,_T_28}; // @[Cat.scala 29:58]
  assign _T_31 = ~ _T_30; // @[convert.scala 21:22]
  assign _T_32 = io_A[2:0]; // @[convert.scala 22:36]
  assign _T_33 = _T_31 < 3'h3; // @[Shift.scala 16:24]
  assign _T_34 = _T_31[1:0]; // @[Shift.scala 17:37]
  assign _T_35 = _T_34[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_32[0:0]; // @[Shift.scala 64:52]
  assign _T_38 = {_T_36,2'h0}; // @[Cat.scala 29:58]
  assign _T_39 = _T_35 ? _T_38 : _T_32; // @[Shift.scala 64:27]
  assign _T_40 = _T_34[0:0]; // @[Shift.scala 66:70]
  assign _T_42 = _T_39[1:0]; // @[Shift.scala 64:52]
  assign _T_43 = {_T_42,1'h0}; // @[Cat.scala 29:58]
  assign _T_44 = _T_40 ? _T_43 : _T_39; // @[Shift.scala 64:27]
  assign decA_fraction = _T_33 ? _T_44 : 3'h0; // @[Shift.scala 16:10]
  assign _T_48 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_50 = _T_3 ? _T_31 : _T_30; // @[convert.scala 25:42]
  assign _T_51 = {_T_48,_T_50}; // @[Cat.scala 29:58]
  assign _T_53 = io_A[4:0]; // @[convert.scala 29:56]
  assign _T_54 = _T_53 != 5'h0; // @[convert.scala 29:60]
  assign _T_55 = ~ _T_54; // @[convert.scala 29:41]
  assign _T_58 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_58 & _T_55; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_51); // @[convert.scala 32:24]
  assign _T_67 = io_B[5]; // @[convert.scala 18:24]
  assign _T_68 = io_B[4]; // @[convert.scala 18:40]
  assign _T_69 = _T_67 ^ _T_68; // @[convert.scala 18:36]
  assign _T_70 = io_B[4:1]; // @[convert.scala 19:24]
  assign _T_71 = io_B[3:0]; // @[convert.scala 19:43]
  assign _T_72 = _T_70 ^ _T_71; // @[convert.scala 19:39]
  assign _T_73 = _T_72[3:2]; // @[LZD.scala 43:32]
  assign _T_74 = _T_73 != 2'h0; // @[LZD.scala 39:14]
  assign _T_75 = _T_73[1]; // @[LZD.scala 39:21]
  assign _T_76 = _T_73[0]; // @[LZD.scala 39:30]
  assign _T_77 = ~ _T_76; // @[LZD.scala 39:27]
  assign _T_78 = _T_75 | _T_77; // @[LZD.scala 39:25]
  assign _T_79 = {_T_74,_T_78}; // @[Cat.scala 29:58]
  assign _T_80 = _T_72[1:0]; // @[LZD.scala 44:32]
  assign _T_81 = _T_80 != 2'h0; // @[LZD.scala 39:14]
  assign _T_82 = _T_80[1]; // @[LZD.scala 39:21]
  assign _T_83 = _T_80[0]; // @[LZD.scala 39:30]
  assign _T_84 = ~ _T_83; // @[LZD.scala 39:27]
  assign _T_85 = _T_82 | _T_84; // @[LZD.scala 39:25]
  assign _T_86 = {_T_81,_T_85}; // @[Cat.scala 29:58]
  assign _T_87 = _T_79[1]; // @[Shift.scala 12:21]
  assign _T_88 = _T_86[1]; // @[Shift.scala 12:21]
  assign _T_89 = _T_87 | _T_88; // @[LZD.scala 49:16]
  assign _T_90 = ~ _T_88; // @[LZD.scala 49:27]
  assign _T_91 = _T_87 | _T_90; // @[LZD.scala 49:25]
  assign _T_92 = _T_79[0:0]; // @[LZD.scala 49:47]
  assign _T_93 = _T_86[0:0]; // @[LZD.scala 49:59]
  assign _T_94 = _T_87 ? _T_92 : _T_93; // @[LZD.scala 49:35]
  assign _T_96 = {_T_89,_T_91,_T_94}; // @[Cat.scala 29:58]
  assign _T_97 = ~ _T_96; // @[convert.scala 21:22]
  assign _T_98 = io_B[2:0]; // @[convert.scala 22:36]
  assign _T_99 = _T_97 < 3'h3; // @[Shift.scala 16:24]
  assign _T_100 = _T_97[1:0]; // @[Shift.scala 17:37]
  assign _T_101 = _T_100[1]; // @[Shift.scala 12:21]
  assign _T_102 = _T_98[0:0]; // @[Shift.scala 64:52]
  assign _T_104 = {_T_102,2'h0}; // @[Cat.scala 29:58]
  assign _T_105 = _T_101 ? _T_104 : _T_98; // @[Shift.scala 64:27]
  assign _T_106 = _T_100[0:0]; // @[Shift.scala 66:70]
  assign _T_108 = _T_105[1:0]; // @[Shift.scala 64:52]
  assign _T_109 = {_T_108,1'h0}; // @[Cat.scala 29:58]
  assign _T_110 = _T_106 ? _T_109 : _T_105; // @[Shift.scala 64:27]
  assign decB_fraction = _T_99 ? _T_110 : 3'h0; // @[Shift.scala 16:10]
  assign _T_114 = _T_69 == 1'h0; // @[convert.scala 25:26]
  assign _T_116 = _T_69 ? _T_97 : _T_96; // @[convert.scala 25:42]
  assign _T_117 = {_T_114,_T_116}; // @[Cat.scala 29:58]
  assign _T_119 = io_B[4:0]; // @[convert.scala 29:56]
  assign _T_120 = _T_119 != 5'h0; // @[convert.scala 29:60]
  assign _T_121 = ~ _T_120; // @[convert.scala 29:41]
  assign _T_124 = _T_67 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_124 & _T_121; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_117); // @[convert.scala 32:24]
  assign aGTb = $signed(decA_scale) > $signed(decB_scale); // @[Sig_op.scala 38:32]
  assign smallerExp = aGTb ? $signed(decB_scale) : $signed(decA_scale); // @[Sig_op.scala 42:24]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[Sig_op.scala 43:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[Sig_op.scala 44:24]
  assign smallerZero = aGTb ? decB_isZero : decA_isZero; // @[Sig_op.scala 45:24]
  assign _T_136 = $signed(io_greaterExp) - $signed(smallerExp); // @[Sig_op.scala 46:35]
  assign scale_diff = $signed(_T_136); // @[Sig_op.scala 46:35]
  assign _T_137 = io_smallerSign | smallerZero; // @[Sig_op.scala 51:53]
  assign _T_138 = ~ _T_137; // @[Sig_op.scala 51:36]
  assign _T_141 = {io_smallerSign,_T_138,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_142 = $unsigned(scale_diff); // @[Sig_op.scala 51:124]
  assign _T_143 = _T_142 < 4'h8; // @[Shift.scala 39:24]
  assign _T_144 = _T_142[2:0]; // @[Shift.scala 40:44]
  assign _T_145 = _T_141[7:4]; // @[Shift.scala 90:30]
  assign _T_146 = _T_141[3:0]; // @[Shift.scala 90:48]
  assign _T_147 = _T_146 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{3'd0}, _T_147}; // @[Shift.scala 90:39]
  assign _T_148 = _T_145 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_149 = _T_144[2]; // @[Shift.scala 12:21]
  assign _T_150 = _T_141[7]; // @[Shift.scala 12:21]
  assign _T_152 = _T_150 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_153 = {_T_152,_T_148}; // @[Cat.scala 29:58]
  assign _T_154 = _T_149 ? _T_153 : _T_141; // @[Shift.scala 91:22]
  assign _T_155 = _T_144[1:0]; // @[Shift.scala 92:77]
  assign _T_156 = _T_154[7:2]; // @[Shift.scala 90:30]
  assign _T_157 = _T_154[1:0]; // @[Shift.scala 90:48]
  assign _T_158 = _T_157 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{5'd0}, _T_158}; // @[Shift.scala 90:39]
  assign _T_159 = _T_156 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_160 = _T_155[1]; // @[Shift.scala 12:21]
  assign _T_161 = _T_154[7]; // @[Shift.scala 12:21]
  assign _T_163 = _T_161 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_164 = {_T_163,_T_159}; // @[Cat.scala 29:58]
  assign _T_165 = _T_160 ? _T_164 : _T_154; // @[Shift.scala 91:22]
  assign _T_166 = _T_155[0:0]; // @[Shift.scala 92:77]
  assign _T_167 = _T_165[7:1]; // @[Shift.scala 90:30]
  assign _T_168 = _T_165[0:0]; // @[Shift.scala 90:48]
  assign _GEN_2 = {{6'd0}, _T_168}; // @[Shift.scala 90:39]
  assign _T_170 = _T_167 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_172 = _T_165[7]; // @[Shift.scala 12:21]
  assign _T_173 = {_T_172,_T_170}; // @[Cat.scala 29:58]
  assign _T_174 = _T_166 ? _T_173 : _T_165; // @[Shift.scala 91:22]
  assign _T_177 = _T_150 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_178 = ~ io_greaterSign; // @[Sig_op.scala 57:40]
  assign _T_179 = {io_greaterSign,_T_178}; // @[Cat.scala 29:58]
  assign io_greaterSign = aGTb ? _T_1 : _T_67; // @[Sig_op.scala 39:18]
  assign io_smallerSign = aGTb ? _T_67 : _T_1; // @[Sig_op.scala 40:18]
  assign io_greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[Sig_op.scala 41:18]
  assign io_greaterSig = {_T_179,greaterFrac}; // @[Sig_op.scala 57:17]
  assign io_smallerSig = _T_143 ? _T_174 : _T_177; // @[Sig_op.scala 52:17]
  assign io_AisNar = _T_1 & _T_55; // @[Sig_op.scala 47:13]
  assign io_BisNar = _T_67 & _T_121; // @[Sig_op.scala 48:13]
  assign io_AisZero = _T_58 & _T_55; // @[Sig_op.scala 49:14]
  assign io_BisZero = _T_124 & _T_121; // @[Sig_op.scala 50:14]
endmodule
