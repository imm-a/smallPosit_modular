module ILZD9(
  input        clock,
  input        reset,
  input  [8:0] io_in,
  output [3:0] io_out
);
  wire [7:0] _T; // @[LZD.scala 43:32]
  wire [3:0] _T_1; // @[LZD.scala 43:32]
  wire [1:0] _T_2; // @[LZD.scala 43:32]
  wire  _T_3; // @[LZD.scala 39:14]
  wire  _T_4; // @[LZD.scala 39:21]
  wire  _T_5; // @[LZD.scala 39:30]
  wire  _T_6; // @[LZD.scala 39:27]
  wire  _T_7; // @[LZD.scala 39:25]
  wire [1:0] _T_8; // @[Cat.scala 29:58]
  wire [1:0] _T_9; // @[LZD.scala 44:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire  _T_16; // @[Shift.scala 12:21]
  wire  _T_17; // @[Shift.scala 12:21]
  wire  _T_18; // @[LZD.scala 49:16]
  wire  _T_19; // @[LZD.scala 49:27]
  wire  _T_20; // @[LZD.scala 49:25]
  wire  _T_21; // @[LZD.scala 49:47]
  wire  _T_22; // @[LZD.scala 49:59]
  wire  _T_23; // @[LZD.scala 49:35]
  wire [2:0] _T_25; // @[Cat.scala 29:58]
  wire [3:0] _T_26; // @[LZD.scala 44:32]
  wire [1:0] _T_27; // @[LZD.scala 43:32]
  wire  _T_28; // @[LZD.scala 39:14]
  wire  _T_29; // @[LZD.scala 39:21]
  wire  _T_30; // @[LZD.scala 39:30]
  wire  _T_31; // @[LZD.scala 39:27]
  wire  _T_32; // @[LZD.scala 39:25]
  wire [1:0] _T_33; // @[Cat.scala 29:58]
  wire [1:0] _T_34; // @[LZD.scala 44:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire  _T_41; // @[Shift.scala 12:21]
  wire  _T_42; // @[Shift.scala 12:21]
  wire  _T_43; // @[LZD.scala 49:16]
  wire  _T_44; // @[LZD.scala 49:27]
  wire  _T_45; // @[LZD.scala 49:25]
  wire  _T_46; // @[LZD.scala 49:47]
  wire  _T_47; // @[LZD.scala 49:59]
  wire  _T_48; // @[LZD.scala 49:35]
  wire [2:0] _T_50; // @[Cat.scala 29:58]
  wire  _T_51; // @[Shift.scala 12:21]
  wire  _T_52; // @[Shift.scala 12:21]
  wire  _T_53; // @[LZD.scala 49:16]
  wire  _T_54; // @[LZD.scala 49:27]
  wire  _T_55; // @[LZD.scala 49:25]
  wire [1:0] _T_56; // @[LZD.scala 49:47]
  wire [1:0] _T_57; // @[LZD.scala 49:59]
  wire [1:0] _T_58; // @[LZD.scala 49:35]
  wire [3:0] _T_60; // @[Cat.scala 29:58]
  wire  _T_61; // @[LZD.scala 44:32]
  wire  _T_63; // @[Shift.scala 12:21]
  wire [2:0] _T_66; // @[Cat.scala 29:58]
  wire [2:0] _T_67; // @[LZD.scala 55:32]
  wire [2:0] _T_68; // @[LZD.scala 55:20]
  assign _T = io_in[8:1]; // @[LZD.scala 43:32]
  assign _T_1 = _T[7:4]; // @[LZD.scala 43:32]
  assign _T_2 = _T_1[3:2]; // @[LZD.scala 43:32]
  assign _T_3 = _T_2 != 2'h0; // @[LZD.scala 39:14]
  assign _T_4 = _T_2[1]; // @[LZD.scala 39:21]
  assign _T_5 = _T_2[0]; // @[LZD.scala 39:30]
  assign _T_6 = ~ _T_5; // @[LZD.scala 39:27]
  assign _T_7 = _T_4 | _T_6; // @[LZD.scala 39:25]
  assign _T_8 = {_T_3,_T_7}; // @[Cat.scala 29:58]
  assign _T_9 = _T_1[1:0]; // @[LZD.scala 44:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1]; // @[Shift.scala 12:21]
  assign _T_17 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_18 = _T_16 | _T_17; // @[LZD.scala 49:16]
  assign _T_19 = ~ _T_17; // @[LZD.scala 49:27]
  assign _T_20 = _T_16 | _T_19; // @[LZD.scala 49:25]
  assign _T_21 = _T_8[0:0]; // @[LZD.scala 49:47]
  assign _T_22 = _T_15[0:0]; // @[LZD.scala 49:59]
  assign _T_23 = _T_16 ? _T_21 : _T_22; // @[LZD.scala 49:35]
  assign _T_25 = {_T_18,_T_20,_T_23}; // @[Cat.scala 29:58]
  assign _T_26 = _T[3:0]; // @[LZD.scala 44:32]
  assign _T_27 = _T_26[3:2]; // @[LZD.scala 43:32]
  assign _T_28 = _T_27 != 2'h0; // @[LZD.scala 39:14]
  assign _T_29 = _T_27[1]; // @[LZD.scala 39:21]
  assign _T_30 = _T_27[0]; // @[LZD.scala 39:30]
  assign _T_31 = ~ _T_30; // @[LZD.scala 39:27]
  assign _T_32 = _T_29 | _T_31; // @[LZD.scala 39:25]
  assign _T_33 = {_T_28,_T_32}; // @[Cat.scala 29:58]
  assign _T_34 = _T_26[1:0]; // @[LZD.scala 44:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1]; // @[Shift.scala 12:21]
  assign _T_42 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_43 = _T_41 | _T_42; // @[LZD.scala 49:16]
  assign _T_44 = ~ _T_42; // @[LZD.scala 49:27]
  assign _T_45 = _T_41 | _T_44; // @[LZD.scala 49:25]
  assign _T_46 = _T_33[0:0]; // @[LZD.scala 49:47]
  assign _T_47 = _T_40[0:0]; // @[LZD.scala 49:59]
  assign _T_48 = _T_41 ? _T_46 : _T_47; // @[LZD.scala 49:35]
  assign _T_50 = {_T_43,_T_45,_T_48}; // @[Cat.scala 29:58]
  assign _T_51 = _T_25[2]; // @[Shift.scala 12:21]
  assign _T_52 = _T_50[2]; // @[Shift.scala 12:21]
  assign _T_53 = _T_51 | _T_52; // @[LZD.scala 49:16]
  assign _T_54 = ~ _T_52; // @[LZD.scala 49:27]
  assign _T_55 = _T_51 | _T_54; // @[LZD.scala 49:25]
  assign _T_56 = _T_25[1:0]; // @[LZD.scala 49:47]
  assign _T_57 = _T_50[1:0]; // @[LZD.scala 49:59]
  assign _T_58 = _T_51 ? _T_56 : _T_57; // @[LZD.scala 49:35]
  assign _T_60 = {_T_53,_T_55,_T_58}; // @[Cat.scala 29:58]
  assign _T_61 = io_in[0:0]; // @[LZD.scala 44:32]
  assign _T_63 = _T_60[3]; // @[Shift.scala 12:21]
  assign _T_66 = {2'h3,_T_61}; // @[Cat.scala 29:58]
  assign _T_67 = _T_60[2:0]; // @[LZD.scala 55:32]
  assign _T_68 = _T_63 ? _T_67 : _T_66; // @[LZD.scala 55:20]
  assign io_out = {_T_63,_T_68}; // @[ILZD.scala 15:10]
endmodule
