module PositFMA7_3(
  input        clock,
  input        reset,
  input        io_inValid,
  input  [1:0] io_fmaOp,
  input  [6:0] io_A,
  input  [6:0] io_B,
  input  [6:0] io_C,
  output [6:0] io_F,
  output       io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [6:0] _T_2; // @[Bitwise.scala 71:12]
  wire [6:0] _T_3; // @[PositFMA.scala 47:41]
  wire [6:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [6:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [6:0] _T_8; // @[Bitwise.scala 71:12]
  wire [6:0] _T_9; // @[PositFMA.scala 48:41]
  wire [6:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [6:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [4:0] _T_16; // @[convert.scala 19:24]
  wire [4:0] _T_17; // @[convert.scala 19:43]
  wire [4:0] _T_18; // @[convert.scala 19:39]
  wire [3:0] _T_19; // @[LZD.scala 43:32]
  wire [1:0] _T_20; // @[LZD.scala 43:32]
  wire  _T_21; // @[LZD.scala 39:14]
  wire  _T_22; // @[LZD.scala 39:21]
  wire  _T_23; // @[LZD.scala 39:30]
  wire  _T_24; // @[LZD.scala 39:27]
  wire  _T_25; // @[LZD.scala 39:25]
  wire [1:0] _T_26; // @[Cat.scala 29:58]
  wire [1:0] _T_27; // @[LZD.scala 44:32]
  wire  _T_28; // @[LZD.scala 39:14]
  wire  _T_29; // @[LZD.scala 39:21]
  wire  _T_30; // @[LZD.scala 39:30]
  wire  _T_31; // @[LZD.scala 39:27]
  wire  _T_32; // @[LZD.scala 39:25]
  wire [1:0] _T_33; // @[Cat.scala 29:58]
  wire  _T_34; // @[Shift.scala 12:21]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[LZD.scala 49:16]
  wire  _T_37; // @[LZD.scala 49:27]
  wire  _T_38; // @[LZD.scala 49:25]
  wire  _T_39; // @[LZD.scala 49:47]
  wire  _T_40; // @[LZD.scala 49:59]
  wire  _T_41; // @[LZD.scala 49:35]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire  _T_44; // @[LZD.scala 44:32]
  wire  _T_46; // @[Shift.scala 12:21]
  wire [1:0] _T_48; // @[Cat.scala 29:58]
  wire [1:0] _T_49; // @[LZD.scala 55:32]
  wire [1:0] _T_50; // @[LZD.scala 55:20]
  wire [2:0] _T_51; // @[Cat.scala 29:58]
  wire [2:0] _T_52; // @[convert.scala 21:22]
  wire [3:0] _T_53; // @[convert.scala 22:36]
  wire  _T_54; // @[Shift.scala 16:24]
  wire [1:0] _T_55; // @[Shift.scala 17:37]
  wire  _T_56; // @[Shift.scala 12:21]
  wire [1:0] _T_57; // @[Shift.scala 64:52]
  wire [3:0] _T_59; // @[Cat.scala 29:58]
  wire [3:0] _T_60; // @[Shift.scala 64:27]
  wire  _T_61; // @[Shift.scala 66:70]
  wire [2:0] _T_63; // @[Shift.scala 64:52]
  wire [3:0] _T_64; // @[Cat.scala 29:58]
  wire [3:0] _T_65; // @[Shift.scala 64:27]
  wire [3:0] _T_66; // @[Shift.scala 16:10]
  wire [2:0] _T_67; // @[convert.scala 23:34]
  wire  decA_fraction; // @[convert.scala 24:34]
  wire  _T_69; // @[convert.scala 25:26]
  wire [2:0] _T_71; // @[convert.scala 25:42]
  wire [2:0] _T_74; // @[convert.scala 26:67]
  wire [2:0] _T_75; // @[convert.scala 26:51]
  wire [6:0] _T_76; // @[Cat.scala 29:58]
  wire [5:0] _T_78; // @[convert.scala 29:56]
  wire  _T_79; // @[convert.scala 29:60]
  wire  _T_80; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_83; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [6:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_92; // @[convert.scala 18:24]
  wire  _T_93; // @[convert.scala 18:40]
  wire  _T_94; // @[convert.scala 18:36]
  wire [4:0] _T_95; // @[convert.scala 19:24]
  wire [4:0] _T_96; // @[convert.scala 19:43]
  wire [4:0] _T_97; // @[convert.scala 19:39]
  wire [3:0] _T_98; // @[LZD.scala 43:32]
  wire [1:0] _T_99; // @[LZD.scala 43:32]
  wire  _T_100; // @[LZD.scala 39:14]
  wire  _T_101; // @[LZD.scala 39:21]
  wire  _T_102; // @[LZD.scala 39:30]
  wire  _T_103; // @[LZD.scala 39:27]
  wire  _T_104; // @[LZD.scala 39:25]
  wire [1:0] _T_105; // @[Cat.scala 29:58]
  wire [1:0] _T_106; // @[LZD.scala 44:32]
  wire  _T_107; // @[LZD.scala 39:14]
  wire  _T_108; // @[LZD.scala 39:21]
  wire  _T_109; // @[LZD.scala 39:30]
  wire  _T_110; // @[LZD.scala 39:27]
  wire  _T_111; // @[LZD.scala 39:25]
  wire [1:0] _T_112; // @[Cat.scala 29:58]
  wire  _T_113; // @[Shift.scala 12:21]
  wire  _T_114; // @[Shift.scala 12:21]
  wire  _T_115; // @[LZD.scala 49:16]
  wire  _T_116; // @[LZD.scala 49:27]
  wire  _T_117; // @[LZD.scala 49:25]
  wire  _T_118; // @[LZD.scala 49:47]
  wire  _T_119; // @[LZD.scala 49:59]
  wire  _T_120; // @[LZD.scala 49:35]
  wire [2:0] _T_122; // @[Cat.scala 29:58]
  wire  _T_123; // @[LZD.scala 44:32]
  wire  _T_125; // @[Shift.scala 12:21]
  wire [1:0] _T_127; // @[Cat.scala 29:58]
  wire [1:0] _T_128; // @[LZD.scala 55:32]
  wire [1:0] _T_129; // @[LZD.scala 55:20]
  wire [2:0] _T_130; // @[Cat.scala 29:58]
  wire [2:0] _T_131; // @[convert.scala 21:22]
  wire [3:0] _T_132; // @[convert.scala 22:36]
  wire  _T_133; // @[Shift.scala 16:24]
  wire [1:0] _T_134; // @[Shift.scala 17:37]
  wire  _T_135; // @[Shift.scala 12:21]
  wire [1:0] _T_136; // @[Shift.scala 64:52]
  wire [3:0] _T_138; // @[Cat.scala 29:58]
  wire [3:0] _T_139; // @[Shift.scala 64:27]
  wire  _T_140; // @[Shift.scala 66:70]
  wire [2:0] _T_142; // @[Shift.scala 64:52]
  wire [3:0] _T_143; // @[Cat.scala 29:58]
  wire [3:0] _T_144; // @[Shift.scala 64:27]
  wire [3:0] _T_145; // @[Shift.scala 16:10]
  wire [2:0] _T_146; // @[convert.scala 23:34]
  wire  decB_fraction; // @[convert.scala 24:34]
  wire  _T_148; // @[convert.scala 25:26]
  wire [2:0] _T_150; // @[convert.scala 25:42]
  wire [2:0] _T_153; // @[convert.scala 26:67]
  wire [2:0] _T_154; // @[convert.scala 26:51]
  wire [6:0] _T_155; // @[Cat.scala 29:58]
  wire [5:0] _T_157; // @[convert.scala 29:56]
  wire  _T_158; // @[convert.scala 29:60]
  wire  _T_159; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_162; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [6:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_171; // @[convert.scala 18:24]
  wire  _T_172; // @[convert.scala 18:40]
  wire  _T_173; // @[convert.scala 18:36]
  wire [4:0] _T_174; // @[convert.scala 19:24]
  wire [4:0] _T_175; // @[convert.scala 19:43]
  wire [4:0] _T_176; // @[convert.scala 19:39]
  wire [3:0] _T_177; // @[LZD.scala 43:32]
  wire [1:0] _T_178; // @[LZD.scala 43:32]
  wire  _T_179; // @[LZD.scala 39:14]
  wire  _T_180; // @[LZD.scala 39:21]
  wire  _T_181; // @[LZD.scala 39:30]
  wire  _T_182; // @[LZD.scala 39:27]
  wire  _T_183; // @[LZD.scala 39:25]
  wire [1:0] _T_184; // @[Cat.scala 29:58]
  wire [1:0] _T_185; // @[LZD.scala 44:32]
  wire  _T_186; // @[LZD.scala 39:14]
  wire  _T_187; // @[LZD.scala 39:21]
  wire  _T_188; // @[LZD.scala 39:30]
  wire  _T_189; // @[LZD.scala 39:27]
  wire  _T_190; // @[LZD.scala 39:25]
  wire [1:0] _T_191; // @[Cat.scala 29:58]
  wire  _T_192; // @[Shift.scala 12:21]
  wire  _T_193; // @[Shift.scala 12:21]
  wire  _T_194; // @[LZD.scala 49:16]
  wire  _T_195; // @[LZD.scala 49:27]
  wire  _T_196; // @[LZD.scala 49:25]
  wire  _T_197; // @[LZD.scala 49:47]
  wire  _T_198; // @[LZD.scala 49:59]
  wire  _T_199; // @[LZD.scala 49:35]
  wire [2:0] _T_201; // @[Cat.scala 29:58]
  wire  _T_202; // @[LZD.scala 44:32]
  wire  _T_204; // @[Shift.scala 12:21]
  wire [1:0] _T_206; // @[Cat.scala 29:58]
  wire [1:0] _T_207; // @[LZD.scala 55:32]
  wire [1:0] _T_208; // @[LZD.scala 55:20]
  wire [2:0] _T_209; // @[Cat.scala 29:58]
  wire [2:0] _T_210; // @[convert.scala 21:22]
  wire [3:0] _T_211; // @[convert.scala 22:36]
  wire  _T_212; // @[Shift.scala 16:24]
  wire [1:0] _T_213; // @[Shift.scala 17:37]
  wire  _T_214; // @[Shift.scala 12:21]
  wire [1:0] _T_215; // @[Shift.scala 64:52]
  wire [3:0] _T_217; // @[Cat.scala 29:58]
  wire [3:0] _T_218; // @[Shift.scala 64:27]
  wire  _T_219; // @[Shift.scala 66:70]
  wire [2:0] _T_221; // @[Shift.scala 64:52]
  wire [3:0] _T_222; // @[Cat.scala 29:58]
  wire [3:0] _T_223; // @[Shift.scala 64:27]
  wire [3:0] _T_224; // @[Shift.scala 16:10]
  wire [2:0] _T_225; // @[convert.scala 23:34]
  wire  decC_fraction; // @[convert.scala 24:34]
  wire  _T_227; // @[convert.scala 25:26]
  wire [2:0] _T_229; // @[convert.scala 25:42]
  wire [2:0] _T_232; // @[convert.scala 26:67]
  wire [2:0] _T_233; // @[convert.scala 26:51]
  wire [6:0] _T_234; // @[Cat.scala 29:58]
  wire [5:0] _T_236; // @[convert.scala 29:56]
  wire  _T_237; // @[convert.scala 29:60]
  wire  _T_238; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_241; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [6:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_249; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_250; // @[PositFMA.scala 59:34]
  wire  _T_251; // @[PositFMA.scala 59:47]
  wire  _T_252; // @[PositFMA.scala 59:45]
  wire [2:0] _T_254; // @[Cat.scala 29:58]
  wire [2:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_255; // @[PositFMA.scala 60:34]
  wire  _T_256; // @[PositFMA.scala 60:47]
  wire  _T_257; // @[PositFMA.scala 60:45]
  wire [2:0] _T_259; // @[Cat.scala 29:58]
  wire [2:0] sigB; // @[PositFMA.scala 60:76]
  wire [5:0] _T_260; // @[PositFMA.scala 62:25]
  wire [5:0] sigP; // @[PositFMA.scala 62:33]
  wire [1:0] head2; // @[PositFMA.scala 63:28]
  wire  _T_261; // @[PositFMA.scala 64:31]
  wire  _T_262; // @[PositFMA.scala 64:25]
  wire  _T_263; // @[PositFMA.scala 64:42]
  wire  addTwo; // @[PositFMA.scala 64:35]
  wire  _T_264; // @[PositFMA.scala 66:23]
  wire  _T_265; // @[PositFMA.scala 66:49]
  wire  addOne; // @[PositFMA.scala 66:43]
  wire [1:0] _T_266; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 67:39]
  wire  mulSign; // @[PositFMA.scala 68:28]
  wire [7:0] _T_267; // @[PositFMA.scala 70:30]
  wire [7:0] _GEN_12; // @[PositFMA.scala 70:44]
  wire [7:0] _T_269; // @[PositFMA.scala 70:44]
  wire [7:0] mulScale; // @[PositFMA.scala 70:44]
  wire [3:0] _T_270; // @[PositFMA.scala 73:29]
  wire [2:0] _T_271; // @[PositFMA.scala 74:29]
  wire [3:0] _T_272; // @[PositFMA.scala 74:48]
  wire [3:0] mulSigTmp; // @[PositFMA.scala 71:22]
  wire  _T_274; // @[PositFMA.scala 78:39]
  wire  _T_275; // @[PositFMA.scala 78:43]
  wire [2:0] _T_276; // @[PositFMA.scala 79:39]
  wire [4:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [4:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [7:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [6:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_302; // @[PositFMA.scala 108:29]
  wire  _T_303; // @[PositFMA.scala 108:47]
  wire  _T_304; // @[PositFMA.scala 108:45]
  wire [4:0] extAddSig; // @[Cat.scala 29:58]
  wire [7:0] _GEN_13; // @[PositFMA.scala 112:39]
  wire  mulGreater; // @[PositFMA.scala 112:39]
  wire [7:0] greaterScale; // @[PositFMA.scala 113:26]
  wire [7:0] smallerScale; // @[PositFMA.scala 114:26]
  wire [7:0] _T_308; // @[PositFMA.scala 115:36]
  wire [7:0] scaleDiff; // @[PositFMA.scala 115:36]
  wire [4:0] greaterSig; // @[PositFMA.scala 116:26]
  wire [4:0] smallerSigTmp; // @[PositFMA.scala 117:26]
  wire [7:0] _T_309; // @[PositFMA.scala 118:69]
  wire  _T_310; // @[Shift.scala 39:24]
  wire [2:0] _T_311; // @[Shift.scala 40:44]
  wire  _T_312; // @[Shift.scala 90:30]
  wire [3:0] _T_313; // @[Shift.scala 90:48]
  wire  _T_314; // @[Shift.scala 90:57]
  wire  _T_315; // @[Shift.scala 90:39]
  wire  _T_316; // @[Shift.scala 12:21]
  wire  _T_317; // @[Shift.scala 12:21]
  wire [3:0] _T_319; // @[Bitwise.scala 71:12]
  wire [4:0] _T_320; // @[Cat.scala 29:58]
  wire [4:0] _T_321; // @[Shift.scala 91:22]
  wire [1:0] _T_322; // @[Shift.scala 92:77]
  wire [2:0] _T_323; // @[Shift.scala 90:30]
  wire [1:0] _T_324; // @[Shift.scala 90:48]
  wire  _T_325; // @[Shift.scala 90:57]
  wire [2:0] _GEN_14; // @[Shift.scala 90:39]
  wire [2:0] _T_326; // @[Shift.scala 90:39]
  wire  _T_327; // @[Shift.scala 12:21]
  wire  _T_328; // @[Shift.scala 12:21]
  wire [1:0] _T_330; // @[Bitwise.scala 71:12]
  wire [4:0] _T_331; // @[Cat.scala 29:58]
  wire [4:0] _T_332; // @[Shift.scala 91:22]
  wire  _T_333; // @[Shift.scala 92:77]
  wire [3:0] _T_334; // @[Shift.scala 90:30]
  wire  _T_335; // @[Shift.scala 90:48]
  wire [3:0] _GEN_15; // @[Shift.scala 90:39]
  wire [3:0] _T_337; // @[Shift.scala 90:39]
  wire  _T_339; // @[Shift.scala 12:21]
  wire [4:0] _T_340; // @[Cat.scala 29:58]
  wire [4:0] _T_341; // @[Shift.scala 91:22]
  wire [4:0] _T_344; // @[Bitwise.scala 71:12]
  wire [4:0] smallerSig; // @[Shift.scala 39:10]
  wire [5:0] rawSumSig; // @[PositFMA.scala 119:34]
  wire  _T_345; // @[PositFMA.scala 120:42]
  wire  _T_346; // @[PositFMA.scala 120:46]
  wire  _T_347; // @[PositFMA.scala 120:79]
  wire  sumSign; // @[PositFMA.scala 120:63]
  wire [4:0] _T_349; // @[PositFMA.scala 121:50]
  wire [5:0] signSumSig; // @[Cat.scala 29:58]
  wire [4:0] _T_350; // @[PositFMA.scala 126:33]
  wire [4:0] _T_351; // @[PositFMA.scala 126:68]
  wire [4:0] sumXor; // @[PositFMA.scala 126:51]
  wire [3:0] _T_352; // @[LZD.scala 43:32]
  wire [1:0] _T_353; // @[LZD.scala 43:32]
  wire  _T_354; // @[LZD.scala 39:14]
  wire  _T_355; // @[LZD.scala 39:21]
  wire  _T_356; // @[LZD.scala 39:30]
  wire  _T_357; // @[LZD.scala 39:27]
  wire  _T_358; // @[LZD.scala 39:25]
  wire [1:0] _T_359; // @[Cat.scala 29:58]
  wire [1:0] _T_360; // @[LZD.scala 44:32]
  wire  _T_361; // @[LZD.scala 39:14]
  wire  _T_362; // @[LZD.scala 39:21]
  wire  _T_363; // @[LZD.scala 39:30]
  wire  _T_364; // @[LZD.scala 39:27]
  wire  _T_365; // @[LZD.scala 39:25]
  wire [1:0] _T_366; // @[Cat.scala 29:58]
  wire  _T_367; // @[Shift.scala 12:21]
  wire  _T_368; // @[Shift.scala 12:21]
  wire  _T_369; // @[LZD.scala 49:16]
  wire  _T_370; // @[LZD.scala 49:27]
  wire  _T_371; // @[LZD.scala 49:25]
  wire  _T_372; // @[LZD.scala 49:47]
  wire  _T_373; // @[LZD.scala 49:59]
  wire  _T_374; // @[LZD.scala 49:35]
  wire [2:0] _T_376; // @[Cat.scala 29:58]
  wire  _T_377; // @[LZD.scala 44:32]
  wire  _T_379; // @[Shift.scala 12:21]
  wire [1:0] _T_381; // @[Cat.scala 29:58]
  wire [1:0] _T_382; // @[LZD.scala 55:32]
  wire [1:0] _T_383; // @[LZD.scala 55:20]
  wire [2:0] sumLZD; // @[Cat.scala 29:58]
  wire [2:0] shiftValue; // @[PositFMA.scala 128:24]
  wire [3:0] _T_384; // @[PositFMA.scala 129:38]
  wire  _T_385; // @[Shift.scala 16:24]
  wire [1:0] _T_386; // @[Shift.scala 17:37]
  wire  _T_387; // @[Shift.scala 12:21]
  wire [1:0] _T_388; // @[Shift.scala 64:52]
  wire [3:0] _T_390; // @[Cat.scala 29:58]
  wire [3:0] _T_391; // @[Shift.scala 64:27]
  wire  _T_392; // @[Shift.scala 66:70]
  wire [2:0] _T_394; // @[Shift.scala 64:52]
  wire [3:0] _T_395; // @[Cat.scala 29:58]
  wire [3:0] _T_396; // @[Shift.scala 64:27]
  wire [3:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [7:0] _T_398; // @[PositFMA.scala 132:36]
  wire [7:0] _T_399; // @[PositFMA.scala 132:36]
  wire [3:0] _T_400; // @[Cat.scala 29:58]
  wire [3:0] _T_401; // @[PositFMA.scala 132:61]
  wire [7:0] _GEN_16; // @[PositFMA.scala 132:42]
  wire [7:0] _T_403; // @[PositFMA.scala 132:42]
  wire [7:0] sumScale; // @[PositFMA.scala 132:42]
  wire  sumFrac; // @[PositFMA.scala 133:41]
  wire [2:0] grsTmp; // @[PositFMA.scala 136:41]
  wire [1:0] _T_404; // @[PositFMA.scala 139:40]
  wire  _T_405; // @[PositFMA.scala 139:56]
  wire  underflow; // @[PositFMA.scala 146:32]
  wire  overflow; // @[PositFMA.scala 147:32]
  wire  _T_407; // @[PositFMA.scala 156:32]
  wire  decF_isZero; // @[PositFMA.scala 156:20]
  wire [7:0] _T_409; // @[Mux.scala 87:16]
  wire [7:0] _T_410; // @[Mux.scala 87:16]
  wire [6:0] _GEN_17; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  wire [6:0] decF_scale; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  wire [2:0] _T_411; // @[convert.scala 46:61]
  wire [2:0] _T_412; // @[convert.scala 46:52]
  wire [2:0] _T_414; // @[convert.scala 46:42]
  wire [3:0] _T_415; // @[convert.scala 48:34]
  wire  _T_416; // @[convert.scala 49:36]
  wire [3:0] _T_418; // @[convert.scala 50:36]
  wire [3:0] _T_419; // @[convert.scala 50:36]
  wire [3:0] _T_420; // @[convert.scala 50:28]
  wire  _T_421; // @[convert.scala 51:31]
  wire  _T_422; // @[convert.scala 52:43]
  wire [8:0] _T_426; // @[Cat.scala 29:58]
  wire [3:0] _T_427; // @[Shift.scala 39:17]
  wire  _T_428; // @[Shift.scala 39:24]
  wire  _T_430; // @[Shift.scala 90:30]
  wire [7:0] _T_431; // @[Shift.scala 90:48]
  wire  _T_432; // @[Shift.scala 90:57]
  wire  _T_433; // @[Shift.scala 90:39]
  wire  _T_434; // @[Shift.scala 12:21]
  wire  _T_435; // @[Shift.scala 12:21]
  wire [7:0] _T_437; // @[Bitwise.scala 71:12]
  wire [8:0] _T_438; // @[Cat.scala 29:58]
  wire [8:0] _T_439; // @[Shift.scala 91:22]
  wire [2:0] _T_440; // @[Shift.scala 92:77]
  wire [4:0] _T_441; // @[Shift.scala 90:30]
  wire [3:0] _T_442; // @[Shift.scala 90:48]
  wire  _T_443; // @[Shift.scala 90:57]
  wire [4:0] _GEN_18; // @[Shift.scala 90:39]
  wire [4:0] _T_444; // @[Shift.scala 90:39]
  wire  _T_445; // @[Shift.scala 12:21]
  wire  _T_446; // @[Shift.scala 12:21]
  wire [3:0] _T_448; // @[Bitwise.scala 71:12]
  wire [8:0] _T_449; // @[Cat.scala 29:58]
  wire [8:0] _T_450; // @[Shift.scala 91:22]
  wire [1:0] _T_451; // @[Shift.scala 92:77]
  wire [6:0] _T_452; // @[Shift.scala 90:30]
  wire [1:0] _T_453; // @[Shift.scala 90:48]
  wire  _T_454; // @[Shift.scala 90:57]
  wire [6:0] _GEN_19; // @[Shift.scala 90:39]
  wire [6:0] _T_455; // @[Shift.scala 90:39]
  wire  _T_456; // @[Shift.scala 12:21]
  wire  _T_457; // @[Shift.scala 12:21]
  wire [1:0] _T_459; // @[Bitwise.scala 71:12]
  wire [8:0] _T_460; // @[Cat.scala 29:58]
  wire [8:0] _T_461; // @[Shift.scala 91:22]
  wire  _T_462; // @[Shift.scala 92:77]
  wire [7:0] _T_463; // @[Shift.scala 90:30]
  wire  _T_464; // @[Shift.scala 90:48]
  wire [7:0] _GEN_20; // @[Shift.scala 90:39]
  wire [7:0] _T_466; // @[Shift.scala 90:39]
  wire  _T_468; // @[Shift.scala 12:21]
  wire [8:0] _T_469; // @[Cat.scala 29:58]
  wire [8:0] _T_470; // @[Shift.scala 91:22]
  wire [8:0] _T_473; // @[Bitwise.scala 71:12]
  wire [8:0] _T_474; // @[Shift.scala 39:10]
  wire  _T_475; // @[convert.scala 55:31]
  wire  _T_476; // @[convert.scala 56:31]
  wire  _T_477; // @[convert.scala 57:31]
  wire  _T_478; // @[convert.scala 58:31]
  wire [5:0] _T_479; // @[convert.scala 59:69]
  wire  _T_480; // @[convert.scala 59:81]
  wire  _T_481; // @[convert.scala 59:50]
  wire  _T_483; // @[convert.scala 60:81]
  wire  _T_484; // @[convert.scala 61:44]
  wire  _T_485; // @[convert.scala 61:52]
  wire  _T_486; // @[convert.scala 61:36]
  wire  _T_487; // @[convert.scala 62:63]
  wire  _T_488; // @[convert.scala 62:103]
  wire  _T_489; // @[convert.scala 62:60]
  wire [5:0] _GEN_21; // @[convert.scala 63:56]
  wire [5:0] _T_492; // @[convert.scala 63:56]
  wire [6:0] _T_493; // @[Cat.scala 29:58]
  reg  _T_497; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [6:0] _T_501; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{6'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{6'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[6]; // @[convert.scala 18:24]
  assign _T_14 = realA[5]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[5:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[4:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[4:1]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[3:2]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20 != 2'h0; // @[LZD.scala 39:14]
  assign _T_22 = _T_20[1]; // @[LZD.scala 39:21]
  assign _T_23 = _T_20[0]; // @[LZD.scala 39:30]
  assign _T_24 = ~ _T_23; // @[LZD.scala 39:27]
  assign _T_25 = _T_22 | _T_24; // @[LZD.scala 39:25]
  assign _T_26 = {_T_21,_T_25}; // @[Cat.scala 29:58]
  assign _T_27 = _T_19[1:0]; // @[LZD.scala 44:32]
  assign _T_28 = _T_27 != 2'h0; // @[LZD.scala 39:14]
  assign _T_29 = _T_27[1]; // @[LZD.scala 39:21]
  assign _T_30 = _T_27[0]; // @[LZD.scala 39:30]
  assign _T_31 = ~ _T_30; // @[LZD.scala 39:27]
  assign _T_32 = _T_29 | _T_31; // @[LZD.scala 39:25]
  assign _T_33 = {_T_28,_T_32}; // @[Cat.scala 29:58]
  assign _T_34 = _T_26[1]; // @[Shift.scala 12:21]
  assign _T_35 = _T_33[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_34 | _T_35; // @[LZD.scala 49:16]
  assign _T_37 = ~ _T_35; // @[LZD.scala 49:27]
  assign _T_38 = _T_34 | _T_37; // @[LZD.scala 49:25]
  assign _T_39 = _T_26[0:0]; // @[LZD.scala 49:47]
  assign _T_40 = _T_33[0:0]; // @[LZD.scala 49:59]
  assign _T_41 = _T_34 ? _T_39 : _T_40; // @[LZD.scala 49:35]
  assign _T_43 = {_T_36,_T_38,_T_41}; // @[Cat.scala 29:58]
  assign _T_44 = _T_18[0:0]; // @[LZD.scala 44:32]
  assign _T_46 = _T_43[2]; // @[Shift.scala 12:21]
  assign _T_48 = {1'h1,_T_44}; // @[Cat.scala 29:58]
  assign _T_49 = _T_43[1:0]; // @[LZD.scala 55:32]
  assign _T_50 = _T_46 ? _T_49 : _T_48; // @[LZD.scala 55:20]
  assign _T_51 = {_T_46,_T_50}; // @[Cat.scala 29:58]
  assign _T_52 = ~ _T_51; // @[convert.scala 21:22]
  assign _T_53 = realA[3:0]; // @[convert.scala 22:36]
  assign _T_54 = _T_52 < 3'h4; // @[Shift.scala 16:24]
  assign _T_55 = _T_52[1:0]; // @[Shift.scala 17:37]
  assign _T_56 = _T_55[1]; // @[Shift.scala 12:21]
  assign _T_57 = _T_53[1:0]; // @[Shift.scala 64:52]
  assign _T_59 = {_T_57,2'h0}; // @[Cat.scala 29:58]
  assign _T_60 = _T_56 ? _T_59 : _T_53; // @[Shift.scala 64:27]
  assign _T_61 = _T_55[0:0]; // @[Shift.scala 66:70]
  assign _T_63 = _T_60[2:0]; // @[Shift.scala 64:52]
  assign _T_64 = {_T_63,1'h0}; // @[Cat.scala 29:58]
  assign _T_65 = _T_61 ? _T_64 : _T_60; // @[Shift.scala 64:27]
  assign _T_66 = _T_54 ? _T_65 : 4'h0; // @[Shift.scala 16:10]
  assign _T_67 = _T_66[3:1]; // @[convert.scala 23:34]
  assign decA_fraction = _T_66[0:0]; // @[convert.scala 24:34]
  assign _T_69 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_71 = _T_15 ? _T_52 : _T_51; // @[convert.scala 25:42]
  assign _T_74 = ~ _T_67; // @[convert.scala 26:67]
  assign _T_75 = _T_13 ? _T_74 : _T_67; // @[convert.scala 26:51]
  assign _T_76 = {_T_69,_T_71,_T_75}; // @[Cat.scala 29:58]
  assign _T_78 = realA[5:0]; // @[convert.scala 29:56]
  assign _T_79 = _T_78 != 6'h0; // @[convert.scala 29:60]
  assign _T_80 = ~ _T_79; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_80; // @[convert.scala 29:39]
  assign _T_83 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_83 & _T_80; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_76); // @[convert.scala 32:24]
  assign _T_92 = io_B[6]; // @[convert.scala 18:24]
  assign _T_93 = io_B[5]; // @[convert.scala 18:40]
  assign _T_94 = _T_92 ^ _T_93; // @[convert.scala 18:36]
  assign _T_95 = io_B[5:1]; // @[convert.scala 19:24]
  assign _T_96 = io_B[4:0]; // @[convert.scala 19:43]
  assign _T_97 = _T_95 ^ _T_96; // @[convert.scala 19:39]
  assign _T_98 = _T_97[4:1]; // @[LZD.scala 43:32]
  assign _T_99 = _T_98[3:2]; // @[LZD.scala 43:32]
  assign _T_100 = _T_99 != 2'h0; // @[LZD.scala 39:14]
  assign _T_101 = _T_99[1]; // @[LZD.scala 39:21]
  assign _T_102 = _T_99[0]; // @[LZD.scala 39:30]
  assign _T_103 = ~ _T_102; // @[LZD.scala 39:27]
  assign _T_104 = _T_101 | _T_103; // @[LZD.scala 39:25]
  assign _T_105 = {_T_100,_T_104}; // @[Cat.scala 29:58]
  assign _T_106 = _T_98[1:0]; // @[LZD.scala 44:32]
  assign _T_107 = _T_106 != 2'h0; // @[LZD.scala 39:14]
  assign _T_108 = _T_106[1]; // @[LZD.scala 39:21]
  assign _T_109 = _T_106[0]; // @[LZD.scala 39:30]
  assign _T_110 = ~ _T_109; // @[LZD.scala 39:27]
  assign _T_111 = _T_108 | _T_110; // @[LZD.scala 39:25]
  assign _T_112 = {_T_107,_T_111}; // @[Cat.scala 29:58]
  assign _T_113 = _T_105[1]; // @[Shift.scala 12:21]
  assign _T_114 = _T_112[1]; // @[Shift.scala 12:21]
  assign _T_115 = _T_113 | _T_114; // @[LZD.scala 49:16]
  assign _T_116 = ~ _T_114; // @[LZD.scala 49:27]
  assign _T_117 = _T_113 | _T_116; // @[LZD.scala 49:25]
  assign _T_118 = _T_105[0:0]; // @[LZD.scala 49:47]
  assign _T_119 = _T_112[0:0]; // @[LZD.scala 49:59]
  assign _T_120 = _T_113 ? _T_118 : _T_119; // @[LZD.scala 49:35]
  assign _T_122 = {_T_115,_T_117,_T_120}; // @[Cat.scala 29:58]
  assign _T_123 = _T_97[0:0]; // @[LZD.scala 44:32]
  assign _T_125 = _T_122[2]; // @[Shift.scala 12:21]
  assign _T_127 = {1'h1,_T_123}; // @[Cat.scala 29:58]
  assign _T_128 = _T_122[1:0]; // @[LZD.scala 55:32]
  assign _T_129 = _T_125 ? _T_128 : _T_127; // @[LZD.scala 55:20]
  assign _T_130 = {_T_125,_T_129}; // @[Cat.scala 29:58]
  assign _T_131 = ~ _T_130; // @[convert.scala 21:22]
  assign _T_132 = io_B[3:0]; // @[convert.scala 22:36]
  assign _T_133 = _T_131 < 3'h4; // @[Shift.scala 16:24]
  assign _T_134 = _T_131[1:0]; // @[Shift.scala 17:37]
  assign _T_135 = _T_134[1]; // @[Shift.scala 12:21]
  assign _T_136 = _T_132[1:0]; // @[Shift.scala 64:52]
  assign _T_138 = {_T_136,2'h0}; // @[Cat.scala 29:58]
  assign _T_139 = _T_135 ? _T_138 : _T_132; // @[Shift.scala 64:27]
  assign _T_140 = _T_134[0:0]; // @[Shift.scala 66:70]
  assign _T_142 = _T_139[2:0]; // @[Shift.scala 64:52]
  assign _T_143 = {_T_142,1'h0}; // @[Cat.scala 29:58]
  assign _T_144 = _T_140 ? _T_143 : _T_139; // @[Shift.scala 64:27]
  assign _T_145 = _T_133 ? _T_144 : 4'h0; // @[Shift.scala 16:10]
  assign _T_146 = _T_145[3:1]; // @[convert.scala 23:34]
  assign decB_fraction = _T_145[0:0]; // @[convert.scala 24:34]
  assign _T_148 = _T_94 == 1'h0; // @[convert.scala 25:26]
  assign _T_150 = _T_94 ? _T_131 : _T_130; // @[convert.scala 25:42]
  assign _T_153 = ~ _T_146; // @[convert.scala 26:67]
  assign _T_154 = _T_92 ? _T_153 : _T_146; // @[convert.scala 26:51]
  assign _T_155 = {_T_148,_T_150,_T_154}; // @[Cat.scala 29:58]
  assign _T_157 = io_B[5:0]; // @[convert.scala 29:56]
  assign _T_158 = _T_157 != 6'h0; // @[convert.scala 29:60]
  assign _T_159 = ~ _T_158; // @[convert.scala 29:41]
  assign decB_isNaR = _T_92 & _T_159; // @[convert.scala 29:39]
  assign _T_162 = _T_92 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_162 & _T_159; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_155); // @[convert.scala 32:24]
  assign _T_171 = realC[6]; // @[convert.scala 18:24]
  assign _T_172 = realC[5]; // @[convert.scala 18:40]
  assign _T_173 = _T_171 ^ _T_172; // @[convert.scala 18:36]
  assign _T_174 = realC[5:1]; // @[convert.scala 19:24]
  assign _T_175 = realC[4:0]; // @[convert.scala 19:43]
  assign _T_176 = _T_174 ^ _T_175; // @[convert.scala 19:39]
  assign _T_177 = _T_176[4:1]; // @[LZD.scala 43:32]
  assign _T_178 = _T_177[3:2]; // @[LZD.scala 43:32]
  assign _T_179 = _T_178 != 2'h0; // @[LZD.scala 39:14]
  assign _T_180 = _T_178[1]; // @[LZD.scala 39:21]
  assign _T_181 = _T_178[0]; // @[LZD.scala 39:30]
  assign _T_182 = ~ _T_181; // @[LZD.scala 39:27]
  assign _T_183 = _T_180 | _T_182; // @[LZD.scala 39:25]
  assign _T_184 = {_T_179,_T_183}; // @[Cat.scala 29:58]
  assign _T_185 = _T_177[1:0]; // @[LZD.scala 44:32]
  assign _T_186 = _T_185 != 2'h0; // @[LZD.scala 39:14]
  assign _T_187 = _T_185[1]; // @[LZD.scala 39:21]
  assign _T_188 = _T_185[0]; // @[LZD.scala 39:30]
  assign _T_189 = ~ _T_188; // @[LZD.scala 39:27]
  assign _T_190 = _T_187 | _T_189; // @[LZD.scala 39:25]
  assign _T_191 = {_T_186,_T_190}; // @[Cat.scala 29:58]
  assign _T_192 = _T_184[1]; // @[Shift.scala 12:21]
  assign _T_193 = _T_191[1]; // @[Shift.scala 12:21]
  assign _T_194 = _T_192 | _T_193; // @[LZD.scala 49:16]
  assign _T_195 = ~ _T_193; // @[LZD.scala 49:27]
  assign _T_196 = _T_192 | _T_195; // @[LZD.scala 49:25]
  assign _T_197 = _T_184[0:0]; // @[LZD.scala 49:47]
  assign _T_198 = _T_191[0:0]; // @[LZD.scala 49:59]
  assign _T_199 = _T_192 ? _T_197 : _T_198; // @[LZD.scala 49:35]
  assign _T_201 = {_T_194,_T_196,_T_199}; // @[Cat.scala 29:58]
  assign _T_202 = _T_176[0:0]; // @[LZD.scala 44:32]
  assign _T_204 = _T_201[2]; // @[Shift.scala 12:21]
  assign _T_206 = {1'h1,_T_202}; // @[Cat.scala 29:58]
  assign _T_207 = _T_201[1:0]; // @[LZD.scala 55:32]
  assign _T_208 = _T_204 ? _T_207 : _T_206; // @[LZD.scala 55:20]
  assign _T_209 = {_T_204,_T_208}; // @[Cat.scala 29:58]
  assign _T_210 = ~ _T_209; // @[convert.scala 21:22]
  assign _T_211 = realC[3:0]; // @[convert.scala 22:36]
  assign _T_212 = _T_210 < 3'h4; // @[Shift.scala 16:24]
  assign _T_213 = _T_210[1:0]; // @[Shift.scala 17:37]
  assign _T_214 = _T_213[1]; // @[Shift.scala 12:21]
  assign _T_215 = _T_211[1:0]; // @[Shift.scala 64:52]
  assign _T_217 = {_T_215,2'h0}; // @[Cat.scala 29:58]
  assign _T_218 = _T_214 ? _T_217 : _T_211; // @[Shift.scala 64:27]
  assign _T_219 = _T_213[0:0]; // @[Shift.scala 66:70]
  assign _T_221 = _T_218[2:0]; // @[Shift.scala 64:52]
  assign _T_222 = {_T_221,1'h0}; // @[Cat.scala 29:58]
  assign _T_223 = _T_219 ? _T_222 : _T_218; // @[Shift.scala 64:27]
  assign _T_224 = _T_212 ? _T_223 : 4'h0; // @[Shift.scala 16:10]
  assign _T_225 = _T_224[3:1]; // @[convert.scala 23:34]
  assign decC_fraction = _T_224[0:0]; // @[convert.scala 24:34]
  assign _T_227 = _T_173 == 1'h0; // @[convert.scala 25:26]
  assign _T_229 = _T_173 ? _T_210 : _T_209; // @[convert.scala 25:42]
  assign _T_232 = ~ _T_225; // @[convert.scala 26:67]
  assign _T_233 = _T_171 ? _T_232 : _T_225; // @[convert.scala 26:51]
  assign _T_234 = {_T_227,_T_229,_T_233}; // @[Cat.scala 29:58]
  assign _T_236 = realC[5:0]; // @[convert.scala 29:56]
  assign _T_237 = _T_236 != 6'h0; // @[convert.scala 29:60]
  assign _T_238 = ~ _T_237; // @[convert.scala 29:41]
  assign decC_isNaR = _T_171 & _T_238; // @[convert.scala 29:39]
  assign _T_241 = _T_171 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_241 & _T_238; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_234); // @[convert.scala 32:24]
  assign _T_249 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_249 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_250 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_251 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_252 = _T_250 & _T_251; // @[PositFMA.scala 59:45]
  assign _T_254 = {_T_13,_T_252,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_254); // @[PositFMA.scala 59:76]
  assign _T_255 = ~ _T_92; // @[PositFMA.scala 60:34]
  assign _T_256 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_257 = _T_255 & _T_256; // @[PositFMA.scala 60:45]
  assign _T_259 = {_T_92,_T_257,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_259); // @[PositFMA.scala 60:76]
  assign _T_260 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 62:25]
  assign sigP = $unsigned(_T_260); // @[PositFMA.scala 62:33]
  assign head2 = sigP[5:4]; // @[PositFMA.scala 63:28]
  assign _T_261 = head2[1]; // @[PositFMA.scala 64:31]
  assign _T_262 = ~ _T_261; // @[PositFMA.scala 64:25]
  assign _T_263 = head2[0]; // @[PositFMA.scala 64:42]
  assign addTwo = _T_262 & _T_263; // @[PositFMA.scala 64:35]
  assign _T_264 = sigP[5]; // @[PositFMA.scala 66:23]
  assign _T_265 = sigP[3]; // @[PositFMA.scala 66:49]
  assign addOne = _T_264 ^ _T_265; // @[PositFMA.scala 66:43]
  assign _T_266 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_266)}; // @[PositFMA.scala 67:39]
  assign mulSign = sigP[5:5]; // @[PositFMA.scala 68:28]
  assign _T_267 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 70:30]
  assign _GEN_12 = {{5{expBias[2]}},expBias}; // @[PositFMA.scala 70:44]
  assign _T_269 = $signed(_T_267) + $signed(_GEN_12); // @[PositFMA.scala 70:44]
  assign mulScale = $signed(_T_269); // @[PositFMA.scala 70:44]
  assign _T_270 = sigP[3:0]; // @[PositFMA.scala 73:29]
  assign _T_271 = sigP[2:0]; // @[PositFMA.scala 74:29]
  assign _T_272 = {_T_271, 1'h0}; // @[PositFMA.scala 74:48]
  assign mulSigTmp = addOne ? _T_270 : _T_272; // @[PositFMA.scala 71:22]
  assign _T_274 = mulSigTmp[3:3]; // @[PositFMA.scala 78:39]
  assign _T_275 = _T_274 | addTwo; // @[PositFMA.scala 78:43]
  assign _T_276 = mulSigTmp[2:0]; // @[PositFMA.scala 79:39]
  assign mulSig = {mulSign,_T_275,_T_276}; // @[Cat.scala 29:58]
  assign _T_302 = ~ addSign_phase2; // @[PositFMA.scala 108:29]
  assign _T_303 = ~ addZero_phase2; // @[PositFMA.scala 108:47]
  assign _T_304 = _T_302 & _T_303; // @[PositFMA.scala 108:45]
  assign extAddSig = {addSign_phase2,_T_304,addFrac_phase2,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[6]}},addScale_phase2}; // @[PositFMA.scala 112:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 112:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[6]}},addScale_phase2}); // @[PositFMA.scala 113:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[6]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 114:26]
  assign _T_308 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 115:36]
  assign scaleDiff = $signed(_T_308); // @[PositFMA.scala 115:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 116:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 117:26]
  assign _T_309 = $unsigned(scaleDiff); // @[PositFMA.scala 118:69]
  assign _T_310 = _T_309 < 8'h5; // @[Shift.scala 39:24]
  assign _T_311 = _T_309[2:0]; // @[Shift.scala 40:44]
  assign _T_312 = smallerSigTmp[4:4]; // @[Shift.scala 90:30]
  assign _T_313 = smallerSigTmp[3:0]; // @[Shift.scala 90:48]
  assign _T_314 = _T_313 != 4'h0; // @[Shift.scala 90:57]
  assign _T_315 = _T_312 | _T_314; // @[Shift.scala 90:39]
  assign _T_316 = _T_311[2]; // @[Shift.scala 12:21]
  assign _T_317 = smallerSigTmp[4]; // @[Shift.scala 12:21]
  assign _T_319 = _T_317 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_320 = {_T_319,_T_315}; // @[Cat.scala 29:58]
  assign _T_321 = _T_316 ? _T_320 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_322 = _T_311[1:0]; // @[Shift.scala 92:77]
  assign _T_323 = _T_321[4:2]; // @[Shift.scala 90:30]
  assign _T_324 = _T_321[1:0]; // @[Shift.scala 90:48]
  assign _T_325 = _T_324 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{2'd0}, _T_325}; // @[Shift.scala 90:39]
  assign _T_326 = _T_323 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_327 = _T_322[1]; // @[Shift.scala 12:21]
  assign _T_328 = _T_321[4]; // @[Shift.scala 12:21]
  assign _T_330 = _T_328 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_331 = {_T_330,_T_326}; // @[Cat.scala 29:58]
  assign _T_332 = _T_327 ? _T_331 : _T_321; // @[Shift.scala 91:22]
  assign _T_333 = _T_322[0:0]; // @[Shift.scala 92:77]
  assign _T_334 = _T_332[4:1]; // @[Shift.scala 90:30]
  assign _T_335 = _T_332[0:0]; // @[Shift.scala 90:48]
  assign _GEN_15 = {{3'd0}, _T_335}; // @[Shift.scala 90:39]
  assign _T_337 = _T_334 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_339 = _T_332[4]; // @[Shift.scala 12:21]
  assign _T_340 = {_T_339,_T_337}; // @[Cat.scala 29:58]
  assign _T_341 = _T_333 ? _T_340 : _T_332; // @[Shift.scala 91:22]
  assign _T_344 = _T_317 ? 5'h1f : 5'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_310 ? _T_341 : _T_344; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 119:34]
  assign _T_345 = mulSig_phase2[4:4]; // @[PositFMA.scala 120:42]
  assign _T_346 = _T_345 ^ addSign_phase2; // @[PositFMA.scala 120:46]
  assign _T_347 = rawSumSig[5:5]; // @[PositFMA.scala 120:79]
  assign sumSign = _T_346 ^ _T_347; // @[PositFMA.scala 120:63]
  assign _T_349 = greaterSig + smallerSig; // @[PositFMA.scala 121:50]
  assign signSumSig = {sumSign,_T_349}; // @[Cat.scala 29:58]
  assign _T_350 = signSumSig[5:1]; // @[PositFMA.scala 126:33]
  assign _T_351 = signSumSig[4:0]; // @[PositFMA.scala 126:68]
  assign sumXor = _T_350 ^ _T_351; // @[PositFMA.scala 126:51]
  assign _T_352 = sumXor[4:1]; // @[LZD.scala 43:32]
  assign _T_353 = _T_352[3:2]; // @[LZD.scala 43:32]
  assign _T_354 = _T_353 != 2'h0; // @[LZD.scala 39:14]
  assign _T_355 = _T_353[1]; // @[LZD.scala 39:21]
  assign _T_356 = _T_353[0]; // @[LZD.scala 39:30]
  assign _T_357 = ~ _T_356; // @[LZD.scala 39:27]
  assign _T_358 = _T_355 | _T_357; // @[LZD.scala 39:25]
  assign _T_359 = {_T_354,_T_358}; // @[Cat.scala 29:58]
  assign _T_360 = _T_352[1:0]; // @[LZD.scala 44:32]
  assign _T_361 = _T_360 != 2'h0; // @[LZD.scala 39:14]
  assign _T_362 = _T_360[1]; // @[LZD.scala 39:21]
  assign _T_363 = _T_360[0]; // @[LZD.scala 39:30]
  assign _T_364 = ~ _T_363; // @[LZD.scala 39:27]
  assign _T_365 = _T_362 | _T_364; // @[LZD.scala 39:25]
  assign _T_366 = {_T_361,_T_365}; // @[Cat.scala 29:58]
  assign _T_367 = _T_359[1]; // @[Shift.scala 12:21]
  assign _T_368 = _T_366[1]; // @[Shift.scala 12:21]
  assign _T_369 = _T_367 | _T_368; // @[LZD.scala 49:16]
  assign _T_370 = ~ _T_368; // @[LZD.scala 49:27]
  assign _T_371 = _T_367 | _T_370; // @[LZD.scala 49:25]
  assign _T_372 = _T_359[0:0]; // @[LZD.scala 49:47]
  assign _T_373 = _T_366[0:0]; // @[LZD.scala 49:59]
  assign _T_374 = _T_367 ? _T_372 : _T_373; // @[LZD.scala 49:35]
  assign _T_376 = {_T_369,_T_371,_T_374}; // @[Cat.scala 29:58]
  assign _T_377 = sumXor[0:0]; // @[LZD.scala 44:32]
  assign _T_379 = _T_376[2]; // @[Shift.scala 12:21]
  assign _T_381 = {1'h1,_T_377}; // @[Cat.scala 29:58]
  assign _T_382 = _T_376[1:0]; // @[LZD.scala 55:32]
  assign _T_383 = _T_379 ? _T_382 : _T_381; // @[LZD.scala 55:20]
  assign sumLZD = {_T_379,_T_383}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 128:24]
  assign _T_384 = signSumSig[3:0]; // @[PositFMA.scala 129:38]
  assign _T_385 = shiftValue < 3'h4; // @[Shift.scala 16:24]
  assign _T_386 = shiftValue[1:0]; // @[Shift.scala 17:37]
  assign _T_387 = _T_386[1]; // @[Shift.scala 12:21]
  assign _T_388 = _T_384[1:0]; // @[Shift.scala 64:52]
  assign _T_390 = {_T_388,2'h0}; // @[Cat.scala 29:58]
  assign _T_391 = _T_387 ? _T_390 : _T_384; // @[Shift.scala 64:27]
  assign _T_392 = _T_386[0:0]; // @[Shift.scala 66:70]
  assign _T_394 = _T_391[2:0]; // @[Shift.scala 64:52]
  assign _T_395 = {_T_394,1'h0}; // @[Cat.scala 29:58]
  assign _T_396 = _T_392 ? _T_395 : _T_391; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_385 ? _T_396 : 4'h0; // @[Shift.scala 16:10]
  assign _T_398 = $signed(greaterScale) + $signed(8'sh2); // @[PositFMA.scala 132:36]
  assign _T_399 = $signed(_T_398); // @[PositFMA.scala 132:36]
  assign _T_400 = {1'h1,_T_379,_T_383}; // @[Cat.scala 29:58]
  assign _T_401 = $signed(_T_400); // @[PositFMA.scala 132:61]
  assign _GEN_16 = {{4{_T_401[3]}},_T_401}; // @[PositFMA.scala 132:42]
  assign _T_403 = $signed(_T_399) + $signed(_GEN_16); // @[PositFMA.scala 132:42]
  assign sumScale = $signed(_T_403); // @[PositFMA.scala 132:42]
  assign sumFrac = normalFracTmp[3:3]; // @[PositFMA.scala 133:41]
  assign grsTmp = normalFracTmp[2:0]; // @[PositFMA.scala 136:41]
  assign _T_404 = grsTmp[2:1]; // @[PositFMA.scala 139:40]
  assign _T_405 = grsTmp[0:0]; // @[PositFMA.scala 139:56]
  assign underflow = $signed(sumScale) < $signed(-8'sh29); // @[PositFMA.scala 146:32]
  assign overflow = $signed(sumScale) > $signed(8'sh28); // @[PositFMA.scala 147:32]
  assign _T_407 = signSumSig != 6'h0; // @[PositFMA.scala 156:32]
  assign decF_isZero = ~ _T_407; // @[PositFMA.scala 156:20]
  assign _T_409 = underflow ? $signed(-8'sh29) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_410 = overflow ? $signed(8'sh28) : $signed(_T_409); // @[Mux.scala 87:16]
  assign _GEN_17 = _T_410[6:0]; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  assign decF_scale = $signed(_GEN_17); // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  assign _T_411 = decF_scale[2:0]; // @[convert.scala 46:61]
  assign _T_412 = ~ _T_411; // @[convert.scala 46:52]
  assign _T_414 = sumSign ? _T_412 : _T_411; // @[convert.scala 46:42]
  assign _T_415 = decF_scale[6:3]; // @[convert.scala 48:34]
  assign _T_416 = _T_415[3:3]; // @[convert.scala 49:36]
  assign _T_418 = ~ _T_415; // @[convert.scala 50:36]
  assign _T_419 = $signed(_T_418); // @[convert.scala 50:36]
  assign _T_420 = _T_416 ? $signed(_T_419) : $signed(_T_415); // @[convert.scala 50:28]
  assign _T_421 = _T_416 ^ sumSign; // @[convert.scala 51:31]
  assign _T_422 = ~ _T_421; // @[convert.scala 52:43]
  assign _T_426 = {_T_422,_T_421,_T_414,sumFrac,_T_404,_T_405}; // @[Cat.scala 29:58]
  assign _T_427 = $unsigned(_T_420); // @[Shift.scala 39:17]
  assign _T_428 = _T_427 < 4'h9; // @[Shift.scala 39:24]
  assign _T_430 = _T_426[8:8]; // @[Shift.scala 90:30]
  assign _T_431 = _T_426[7:0]; // @[Shift.scala 90:48]
  assign _T_432 = _T_431 != 8'h0; // @[Shift.scala 90:57]
  assign _T_433 = _T_430 | _T_432; // @[Shift.scala 90:39]
  assign _T_434 = _T_427[3]; // @[Shift.scala 12:21]
  assign _T_435 = _T_426[8]; // @[Shift.scala 12:21]
  assign _T_437 = _T_435 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_438 = {_T_437,_T_433}; // @[Cat.scala 29:58]
  assign _T_439 = _T_434 ? _T_438 : _T_426; // @[Shift.scala 91:22]
  assign _T_440 = _T_427[2:0]; // @[Shift.scala 92:77]
  assign _T_441 = _T_439[8:4]; // @[Shift.scala 90:30]
  assign _T_442 = _T_439[3:0]; // @[Shift.scala 90:48]
  assign _T_443 = _T_442 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_18 = {{4'd0}, _T_443}; // @[Shift.scala 90:39]
  assign _T_444 = _T_441 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_445 = _T_440[2]; // @[Shift.scala 12:21]
  assign _T_446 = _T_439[8]; // @[Shift.scala 12:21]
  assign _T_448 = _T_446 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_449 = {_T_448,_T_444}; // @[Cat.scala 29:58]
  assign _T_450 = _T_445 ? _T_449 : _T_439; // @[Shift.scala 91:22]
  assign _T_451 = _T_440[1:0]; // @[Shift.scala 92:77]
  assign _T_452 = _T_450[8:2]; // @[Shift.scala 90:30]
  assign _T_453 = _T_450[1:0]; // @[Shift.scala 90:48]
  assign _T_454 = _T_453 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_19 = {{6'd0}, _T_454}; // @[Shift.scala 90:39]
  assign _T_455 = _T_452 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_456 = _T_451[1]; // @[Shift.scala 12:21]
  assign _T_457 = _T_450[8]; // @[Shift.scala 12:21]
  assign _T_459 = _T_457 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_460 = {_T_459,_T_455}; // @[Cat.scala 29:58]
  assign _T_461 = _T_456 ? _T_460 : _T_450; // @[Shift.scala 91:22]
  assign _T_462 = _T_451[0:0]; // @[Shift.scala 92:77]
  assign _T_463 = _T_461[8:1]; // @[Shift.scala 90:30]
  assign _T_464 = _T_461[0:0]; // @[Shift.scala 90:48]
  assign _GEN_20 = {{7'd0}, _T_464}; // @[Shift.scala 90:39]
  assign _T_466 = _T_463 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_468 = _T_461[8]; // @[Shift.scala 12:21]
  assign _T_469 = {_T_468,_T_466}; // @[Cat.scala 29:58]
  assign _T_470 = _T_462 ? _T_469 : _T_461; // @[Shift.scala 91:22]
  assign _T_473 = _T_435 ? 9'h1ff : 9'h0; // @[Bitwise.scala 71:12]
  assign _T_474 = _T_428 ? _T_470 : _T_473; // @[Shift.scala 39:10]
  assign _T_475 = _T_474[3]; // @[convert.scala 55:31]
  assign _T_476 = _T_474[2]; // @[convert.scala 56:31]
  assign _T_477 = _T_474[1]; // @[convert.scala 57:31]
  assign _T_478 = _T_474[0]; // @[convert.scala 58:31]
  assign _T_479 = _T_474[8:3]; // @[convert.scala 59:69]
  assign _T_480 = _T_479 != 6'h0; // @[convert.scala 59:81]
  assign _T_481 = ~ _T_480; // @[convert.scala 59:50]
  assign _T_483 = _T_479 == 6'h3f; // @[convert.scala 60:81]
  assign _T_484 = _T_475 | _T_477; // @[convert.scala 61:44]
  assign _T_485 = _T_484 | _T_478; // @[convert.scala 61:52]
  assign _T_486 = _T_476 & _T_485; // @[convert.scala 61:36]
  assign _T_487 = ~ _T_483; // @[convert.scala 62:63]
  assign _T_488 = _T_487 & _T_486; // @[convert.scala 62:103]
  assign _T_489 = _T_481 | _T_488; // @[convert.scala 62:60]
  assign _GEN_21 = {{5'd0}, _T_489}; // @[convert.scala 63:56]
  assign _T_492 = _T_479 + _GEN_21; // @[convert.scala 63:56]
  assign _T_493 = {sumSign,_T_492}; // @[Cat.scala 29:58]
  assign io_F = _T_501; // @[PositFMA.scala 176:15]
  assign io_outValid = _T_497; // @[PositFMA.scala 175:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulSig_phase2 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_497 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_501 = _RAND_9[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_171;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_497 <= 1'h0;
    end else begin
      _T_497 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_501 <= 7'h40;
      end else begin
        if (decF_isZero) begin
          _T_501 <= 7'h0;
        end else begin
          _T_501 <= _T_493;
        end
      end
    end
  end
endmodule
