module FMA_Dec4_0(
  input        clock,
  input        reset,
  input  [3:0] io_A,
  input  [3:0] io_B,
  input  [3:0] io_C,
  output [2:0] io_sigA,
  output [2:0] io_sigB,
  output       io_outIsNaR,
  output       io_Csign,
  output       io_CisNar,
  output       io_CisZero,
  output       io_Cfrac,
  output [2:0] io_Ascale,
  output [2:0] io_Bscale,
  output [2:0] io_Cscale
);
  wire [4:0] _T_2; // @[FMA_Dec.scala 38:46]
  wire [3:0] realA; // @[FMA_Dec.scala 38:46]
  wire [4:0] _T_5; // @[FMA_Dec.scala 39:46]
  wire [3:0] realC; // @[FMA_Dec.scala 39:46]
  wire  _T_7; // @[convert.scala 18:24]
  wire  _T_8; // @[convert.scala 18:40]
  wire  _T_9; // @[convert.scala 18:36]
  wire [1:0] _T_10; // @[convert.scala 19:24]
  wire [1:0] _T_11; // @[convert.scala 19:43]
  wire [1:0] _T_12; // @[convert.scala 19:39]
  wire  _T_13; // @[LZD.scala 39:14]
  wire  _T_14; // @[LZD.scala 39:21]
  wire  _T_15; // @[LZD.scala 39:30]
  wire  _T_16; // @[LZD.scala 39:27]
  wire  _T_17; // @[LZD.scala 39:25]
  wire [1:0] _T_18; // @[Cat.scala 29:58]
  wire [1:0] _T_19; // @[convert.scala 21:22]
  wire  _T_20; // @[convert.scala 22:36]
  wire  _T_21; // @[Shift.scala 16:24]
  wire  _T_22; // @[Shift.scala 17:37]
  wire  _T_24; // @[Shift.scala 63:39]
  wire  decA_fraction; // @[Shift.scala 16:10]
  wire  _T_28; // @[convert.scala 25:26]
  wire [1:0] _T_30; // @[convert.scala 25:42]
  wire [2:0] _T_31; // @[Cat.scala 29:58]
  wire [2:0] _T_33; // @[convert.scala 29:56]
  wire  _T_34; // @[convert.scala 29:60]
  wire  _T_35; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_38; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire  _T_47; // @[convert.scala 18:24]
  wire  _T_48; // @[convert.scala 18:40]
  wire  _T_49; // @[convert.scala 18:36]
  wire [1:0] _T_50; // @[convert.scala 19:24]
  wire [1:0] _T_51; // @[convert.scala 19:43]
  wire [1:0] _T_52; // @[convert.scala 19:39]
  wire  _T_53; // @[LZD.scala 39:14]
  wire  _T_54; // @[LZD.scala 39:21]
  wire  _T_55; // @[LZD.scala 39:30]
  wire  _T_56; // @[LZD.scala 39:27]
  wire  _T_57; // @[LZD.scala 39:25]
  wire [1:0] _T_58; // @[Cat.scala 29:58]
  wire [1:0] _T_59; // @[convert.scala 21:22]
  wire  _T_60; // @[convert.scala 22:36]
  wire  _T_61; // @[Shift.scala 16:24]
  wire  _T_62; // @[Shift.scala 17:37]
  wire  _T_64; // @[Shift.scala 63:39]
  wire  decB_fraction; // @[Shift.scala 16:10]
  wire  _T_68; // @[convert.scala 25:26]
  wire [1:0] _T_70; // @[convert.scala 25:42]
  wire [2:0] _T_71; // @[Cat.scala 29:58]
  wire [2:0] _T_73; // @[convert.scala 29:56]
  wire  _T_74; // @[convert.scala 29:60]
  wire  _T_75; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_78; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire  _T_87; // @[convert.scala 18:24]
  wire  _T_88; // @[convert.scala 18:40]
  wire  _T_89; // @[convert.scala 18:36]
  wire [1:0] _T_90; // @[convert.scala 19:24]
  wire [1:0] _T_91; // @[convert.scala 19:43]
  wire [1:0] _T_92; // @[convert.scala 19:39]
  wire  _T_93; // @[LZD.scala 39:14]
  wire  _T_94; // @[LZD.scala 39:21]
  wire  _T_95; // @[LZD.scala 39:30]
  wire  _T_96; // @[LZD.scala 39:27]
  wire  _T_97; // @[LZD.scala 39:25]
  wire [1:0] _T_98; // @[Cat.scala 29:58]
  wire [1:0] _T_99; // @[convert.scala 21:22]
  wire  _T_100; // @[convert.scala 22:36]
  wire  _T_101; // @[Shift.scala 16:24]
  wire  _T_102; // @[Shift.scala 17:37]
  wire  _T_104; // @[Shift.scala 63:39]
  wire  _T_108; // @[convert.scala 25:26]
  wire [1:0] _T_110; // @[convert.scala 25:42]
  wire [2:0] _T_111; // @[Cat.scala 29:58]
  wire [2:0] _T_113; // @[convert.scala 29:56]
  wire  _T_114; // @[convert.scala 29:60]
  wire  _T_115; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_118; // @[convert.scala 30:19]
  wire  _T_126; // @[FMA_Dec.scala 46:30]
  wire  _T_128; // @[FMA_Dec.scala 49:34]
  wire  _T_129; // @[FMA_Dec.scala 49:47]
  wire  _T_130; // @[FMA_Dec.scala 49:45]
  wire [2:0] _T_132; // @[Cat.scala 29:58]
  wire  _T_134; // @[FMA_Dec.scala 50:34]
  wire  _T_135; // @[FMA_Dec.scala 50:47]
  wire  _T_136; // @[FMA_Dec.scala 50:45]
  wire [2:0] _T_138; // @[Cat.scala 29:58]
  assign _T_2 = {{1'd0}, io_A}; // @[FMA_Dec.scala 38:46]
  assign realA = _T_2[3:0]; // @[FMA_Dec.scala 38:46]
  assign _T_5 = {{1'd0}, io_C}; // @[FMA_Dec.scala 39:46]
  assign realC = _T_5[3:0]; // @[FMA_Dec.scala 39:46]
  assign _T_7 = realA[3]; // @[convert.scala 18:24]
  assign _T_8 = realA[2]; // @[convert.scala 18:40]
  assign _T_9 = _T_7 ^ _T_8; // @[convert.scala 18:36]
  assign _T_10 = realA[2:1]; // @[convert.scala 19:24]
  assign _T_11 = realA[1:0]; // @[convert.scala 19:43]
  assign _T_12 = _T_10 ^ _T_11; // @[convert.scala 19:39]
  assign _T_13 = _T_12 != 2'h0; // @[LZD.scala 39:14]
  assign _T_14 = _T_12[1]; // @[LZD.scala 39:21]
  assign _T_15 = _T_12[0]; // @[LZD.scala 39:30]
  assign _T_16 = ~ _T_15; // @[LZD.scala 39:27]
  assign _T_17 = _T_14 | _T_16; // @[LZD.scala 39:25]
  assign _T_18 = {_T_13,_T_17}; // @[Cat.scala 29:58]
  assign _T_19 = ~ _T_18; // @[convert.scala 21:22]
  assign _T_20 = realA[0:0]; // @[convert.scala 22:36]
  assign _T_21 = _T_19 < 2'h1; // @[Shift.scala 16:24]
  assign _T_22 = _T_19[0]; // @[Shift.scala 17:37]
  assign _T_24 = _T_22 ? 1'h0 : _T_20; // @[Shift.scala 63:39]
  assign decA_fraction = _T_21 & _T_24; // @[Shift.scala 16:10]
  assign _T_28 = _T_9 == 1'h0; // @[convert.scala 25:26]
  assign _T_30 = _T_9 ? _T_19 : _T_18; // @[convert.scala 25:42]
  assign _T_31 = {_T_28,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = realA[2:0]; // @[convert.scala 29:56]
  assign _T_34 = _T_33 != 3'h0; // @[convert.scala 29:60]
  assign _T_35 = ~ _T_34; // @[convert.scala 29:41]
  assign decA_isNaR = _T_7 & _T_35; // @[convert.scala 29:39]
  assign _T_38 = _T_7 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_38 & _T_35; // @[convert.scala 30:41]
  assign _T_47 = io_B[3]; // @[convert.scala 18:24]
  assign _T_48 = io_B[2]; // @[convert.scala 18:40]
  assign _T_49 = _T_47 ^ _T_48; // @[convert.scala 18:36]
  assign _T_50 = io_B[2:1]; // @[convert.scala 19:24]
  assign _T_51 = io_B[1:0]; // @[convert.scala 19:43]
  assign _T_52 = _T_50 ^ _T_51; // @[convert.scala 19:39]
  assign _T_53 = _T_52 != 2'h0; // @[LZD.scala 39:14]
  assign _T_54 = _T_52[1]; // @[LZD.scala 39:21]
  assign _T_55 = _T_52[0]; // @[LZD.scala 39:30]
  assign _T_56 = ~ _T_55; // @[LZD.scala 39:27]
  assign _T_57 = _T_54 | _T_56; // @[LZD.scala 39:25]
  assign _T_58 = {_T_53,_T_57}; // @[Cat.scala 29:58]
  assign _T_59 = ~ _T_58; // @[convert.scala 21:22]
  assign _T_60 = io_B[0:0]; // @[convert.scala 22:36]
  assign _T_61 = _T_59 < 2'h1; // @[Shift.scala 16:24]
  assign _T_62 = _T_59[0]; // @[Shift.scala 17:37]
  assign _T_64 = _T_62 ? 1'h0 : _T_60; // @[Shift.scala 63:39]
  assign decB_fraction = _T_61 & _T_64; // @[Shift.scala 16:10]
  assign _T_68 = _T_49 == 1'h0; // @[convert.scala 25:26]
  assign _T_70 = _T_49 ? _T_59 : _T_58; // @[convert.scala 25:42]
  assign _T_71 = {_T_68,_T_70}; // @[Cat.scala 29:58]
  assign _T_73 = io_B[2:0]; // @[convert.scala 29:56]
  assign _T_74 = _T_73 != 3'h0; // @[convert.scala 29:60]
  assign _T_75 = ~ _T_74; // @[convert.scala 29:41]
  assign decB_isNaR = _T_47 & _T_75; // @[convert.scala 29:39]
  assign _T_78 = _T_47 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_78 & _T_75; // @[convert.scala 30:41]
  assign _T_87 = realC[3]; // @[convert.scala 18:24]
  assign _T_88 = realC[2]; // @[convert.scala 18:40]
  assign _T_89 = _T_87 ^ _T_88; // @[convert.scala 18:36]
  assign _T_90 = realC[2:1]; // @[convert.scala 19:24]
  assign _T_91 = realC[1:0]; // @[convert.scala 19:43]
  assign _T_92 = _T_90 ^ _T_91; // @[convert.scala 19:39]
  assign _T_93 = _T_92 != 2'h0; // @[LZD.scala 39:14]
  assign _T_94 = _T_92[1]; // @[LZD.scala 39:21]
  assign _T_95 = _T_92[0]; // @[LZD.scala 39:30]
  assign _T_96 = ~ _T_95; // @[LZD.scala 39:27]
  assign _T_97 = _T_94 | _T_96; // @[LZD.scala 39:25]
  assign _T_98 = {_T_93,_T_97}; // @[Cat.scala 29:58]
  assign _T_99 = ~ _T_98; // @[convert.scala 21:22]
  assign _T_100 = realC[0:0]; // @[convert.scala 22:36]
  assign _T_101 = _T_99 < 2'h1; // @[Shift.scala 16:24]
  assign _T_102 = _T_99[0]; // @[Shift.scala 17:37]
  assign _T_104 = _T_102 ? 1'h0 : _T_100; // @[Shift.scala 63:39]
  assign _T_108 = _T_89 == 1'h0; // @[convert.scala 25:26]
  assign _T_110 = _T_89 ? _T_99 : _T_98; // @[convert.scala 25:42]
  assign _T_111 = {_T_108,_T_110}; // @[Cat.scala 29:58]
  assign _T_113 = realC[2:0]; // @[convert.scala 29:56]
  assign _T_114 = _T_113 != 3'h0; // @[convert.scala 29:60]
  assign _T_115 = ~ _T_114; // @[convert.scala 29:41]
  assign decC_isNaR = _T_87 & _T_115; // @[convert.scala 29:39]
  assign _T_118 = _T_87 == 1'h0; // @[convert.scala 30:19]
  assign _T_126 = decA_isNaR | decB_isNaR; // @[FMA_Dec.scala 46:30]
  assign _T_128 = ~ _T_7; // @[FMA_Dec.scala 49:34]
  assign _T_129 = ~ decA_isZero; // @[FMA_Dec.scala 49:47]
  assign _T_130 = _T_128 & _T_129; // @[FMA_Dec.scala 49:45]
  assign _T_132 = {_T_7,_T_130,decA_fraction}; // @[Cat.scala 29:58]
  assign _T_134 = ~ _T_47; // @[FMA_Dec.scala 50:34]
  assign _T_135 = ~ decB_isZero; // @[FMA_Dec.scala 50:47]
  assign _T_136 = _T_134 & _T_135; // @[FMA_Dec.scala 50:45]
  assign _T_138 = {_T_47,_T_136,decB_fraction}; // @[Cat.scala 29:58]
  assign io_sigA = $signed(_T_132); // @[FMA_Dec.scala 49:16]
  assign io_sigB = $signed(_T_138); // @[FMA_Dec.scala 50:16]
  assign io_outIsNaR = _T_126 | decC_isNaR; // @[FMA_Dec.scala 46:16]
  assign io_Csign = realC[3]; // @[FMA_Dec.scala 55:12]
  assign io_CisNar = _T_87 & _T_115; // @[FMA_Dec.scala 51:17]
  assign io_CisZero = _T_118 & _T_115; // @[FMA_Dec.scala 52:17]
  assign io_Cfrac = _T_101 & _T_104; // @[FMA_Dec.scala 53:17]
  assign io_Ascale = $signed(_T_31); // @[FMA_Dec.scala 47:13]
  assign io_Bscale = $signed(_T_71); // @[FMA_Dec.scala 48:13]
  assign io_Cscale = $signed(_T_111); // @[FMA_Dec.scala 54:16]
endmodule
