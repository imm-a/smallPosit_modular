module PositFMA7_0(
  input        clock,
  input        reset,
  input        io_inValid,
  input  [1:0] io_fmaOp,
  input  [6:0] io_A,
  input  [6:0] io_B,
  input  [6:0] io_C,
  output [6:0] io_F,
  output       io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [6:0] _T_2; // @[Bitwise.scala 71:12]
  wire [6:0] _T_3; // @[PositFMA.scala 47:41]
  wire [6:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [6:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [6:0] _T_8; // @[Bitwise.scala 71:12]
  wire [6:0] _T_9; // @[PositFMA.scala 48:41]
  wire [6:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [6:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [4:0] _T_16; // @[convert.scala 19:24]
  wire [4:0] _T_17; // @[convert.scala 19:43]
  wire [4:0] _T_18; // @[convert.scala 19:39]
  wire [3:0] _T_19; // @[LZD.scala 43:32]
  wire [1:0] _T_20; // @[LZD.scala 43:32]
  wire  _T_21; // @[LZD.scala 39:14]
  wire  _T_22; // @[LZD.scala 39:21]
  wire  _T_23; // @[LZD.scala 39:30]
  wire  _T_24; // @[LZD.scala 39:27]
  wire  _T_25; // @[LZD.scala 39:25]
  wire [1:0] _T_26; // @[Cat.scala 29:58]
  wire [1:0] _T_27; // @[LZD.scala 44:32]
  wire  _T_28; // @[LZD.scala 39:14]
  wire  _T_29; // @[LZD.scala 39:21]
  wire  _T_30; // @[LZD.scala 39:30]
  wire  _T_31; // @[LZD.scala 39:27]
  wire  _T_32; // @[LZD.scala 39:25]
  wire [1:0] _T_33; // @[Cat.scala 29:58]
  wire  _T_34; // @[Shift.scala 12:21]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[LZD.scala 49:16]
  wire  _T_37; // @[LZD.scala 49:27]
  wire  _T_38; // @[LZD.scala 49:25]
  wire  _T_39; // @[LZD.scala 49:47]
  wire  _T_40; // @[LZD.scala 49:59]
  wire  _T_41; // @[LZD.scala 49:35]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire  _T_44; // @[LZD.scala 44:32]
  wire  _T_46; // @[Shift.scala 12:21]
  wire [1:0] _T_48; // @[Cat.scala 29:58]
  wire [1:0] _T_49; // @[LZD.scala 55:32]
  wire [1:0] _T_50; // @[LZD.scala 55:20]
  wire [2:0] _T_51; // @[Cat.scala 29:58]
  wire [2:0] _T_52; // @[convert.scala 21:22]
  wire [3:0] _T_53; // @[convert.scala 22:36]
  wire  _T_54; // @[Shift.scala 16:24]
  wire [1:0] _T_55; // @[Shift.scala 17:37]
  wire  _T_56; // @[Shift.scala 12:21]
  wire [1:0] _T_57; // @[Shift.scala 64:52]
  wire [3:0] _T_59; // @[Cat.scala 29:58]
  wire [3:0] _T_60; // @[Shift.scala 64:27]
  wire  _T_61; // @[Shift.scala 66:70]
  wire [2:0] _T_63; // @[Shift.scala 64:52]
  wire [3:0] _T_64; // @[Cat.scala 29:58]
  wire [3:0] _T_65; // @[Shift.scala 64:27]
  wire [3:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_69; // @[convert.scala 25:26]
  wire [2:0] _T_71; // @[convert.scala 25:42]
  wire [3:0] _T_72; // @[Cat.scala 29:58]
  wire [5:0] _T_74; // @[convert.scala 29:56]
  wire  _T_75; // @[convert.scala 29:60]
  wire  _T_76; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_79; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [3:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_88; // @[convert.scala 18:24]
  wire  _T_89; // @[convert.scala 18:40]
  wire  _T_90; // @[convert.scala 18:36]
  wire [4:0] _T_91; // @[convert.scala 19:24]
  wire [4:0] _T_92; // @[convert.scala 19:43]
  wire [4:0] _T_93; // @[convert.scala 19:39]
  wire [3:0] _T_94; // @[LZD.scala 43:32]
  wire [1:0] _T_95; // @[LZD.scala 43:32]
  wire  _T_96; // @[LZD.scala 39:14]
  wire  _T_97; // @[LZD.scala 39:21]
  wire  _T_98; // @[LZD.scala 39:30]
  wire  _T_99; // @[LZD.scala 39:27]
  wire  _T_100; // @[LZD.scala 39:25]
  wire [1:0] _T_101; // @[Cat.scala 29:58]
  wire [1:0] _T_102; // @[LZD.scala 44:32]
  wire  _T_103; // @[LZD.scala 39:14]
  wire  _T_104; // @[LZD.scala 39:21]
  wire  _T_105; // @[LZD.scala 39:30]
  wire  _T_106; // @[LZD.scala 39:27]
  wire  _T_107; // @[LZD.scala 39:25]
  wire [1:0] _T_108; // @[Cat.scala 29:58]
  wire  _T_109; // @[Shift.scala 12:21]
  wire  _T_110; // @[Shift.scala 12:21]
  wire  _T_111; // @[LZD.scala 49:16]
  wire  _T_112; // @[LZD.scala 49:27]
  wire  _T_113; // @[LZD.scala 49:25]
  wire  _T_114; // @[LZD.scala 49:47]
  wire  _T_115; // @[LZD.scala 49:59]
  wire  _T_116; // @[LZD.scala 49:35]
  wire [2:0] _T_118; // @[Cat.scala 29:58]
  wire  _T_119; // @[LZD.scala 44:32]
  wire  _T_121; // @[Shift.scala 12:21]
  wire [1:0] _T_123; // @[Cat.scala 29:58]
  wire [1:0] _T_124; // @[LZD.scala 55:32]
  wire [1:0] _T_125; // @[LZD.scala 55:20]
  wire [2:0] _T_126; // @[Cat.scala 29:58]
  wire [2:0] _T_127; // @[convert.scala 21:22]
  wire [3:0] _T_128; // @[convert.scala 22:36]
  wire  _T_129; // @[Shift.scala 16:24]
  wire [1:0] _T_130; // @[Shift.scala 17:37]
  wire  _T_131; // @[Shift.scala 12:21]
  wire [1:0] _T_132; // @[Shift.scala 64:52]
  wire [3:0] _T_134; // @[Cat.scala 29:58]
  wire [3:0] _T_135; // @[Shift.scala 64:27]
  wire  _T_136; // @[Shift.scala 66:70]
  wire [2:0] _T_138; // @[Shift.scala 64:52]
  wire [3:0] _T_139; // @[Cat.scala 29:58]
  wire [3:0] _T_140; // @[Shift.scala 64:27]
  wire [3:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_144; // @[convert.scala 25:26]
  wire [2:0] _T_146; // @[convert.scala 25:42]
  wire [3:0] _T_147; // @[Cat.scala 29:58]
  wire [5:0] _T_149; // @[convert.scala 29:56]
  wire  _T_150; // @[convert.scala 29:60]
  wire  _T_151; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_154; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [3:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_163; // @[convert.scala 18:24]
  wire  _T_164; // @[convert.scala 18:40]
  wire  _T_165; // @[convert.scala 18:36]
  wire [4:0] _T_166; // @[convert.scala 19:24]
  wire [4:0] _T_167; // @[convert.scala 19:43]
  wire [4:0] _T_168; // @[convert.scala 19:39]
  wire [3:0] _T_169; // @[LZD.scala 43:32]
  wire [1:0] _T_170; // @[LZD.scala 43:32]
  wire  _T_171; // @[LZD.scala 39:14]
  wire  _T_172; // @[LZD.scala 39:21]
  wire  _T_173; // @[LZD.scala 39:30]
  wire  _T_174; // @[LZD.scala 39:27]
  wire  _T_175; // @[LZD.scala 39:25]
  wire [1:0] _T_176; // @[Cat.scala 29:58]
  wire [1:0] _T_177; // @[LZD.scala 44:32]
  wire  _T_178; // @[LZD.scala 39:14]
  wire  _T_179; // @[LZD.scala 39:21]
  wire  _T_180; // @[LZD.scala 39:30]
  wire  _T_181; // @[LZD.scala 39:27]
  wire  _T_182; // @[LZD.scala 39:25]
  wire [1:0] _T_183; // @[Cat.scala 29:58]
  wire  _T_184; // @[Shift.scala 12:21]
  wire  _T_185; // @[Shift.scala 12:21]
  wire  _T_186; // @[LZD.scala 49:16]
  wire  _T_187; // @[LZD.scala 49:27]
  wire  _T_188; // @[LZD.scala 49:25]
  wire  _T_189; // @[LZD.scala 49:47]
  wire  _T_190; // @[LZD.scala 49:59]
  wire  _T_191; // @[LZD.scala 49:35]
  wire [2:0] _T_193; // @[Cat.scala 29:58]
  wire  _T_194; // @[LZD.scala 44:32]
  wire  _T_196; // @[Shift.scala 12:21]
  wire [1:0] _T_198; // @[Cat.scala 29:58]
  wire [1:0] _T_199; // @[LZD.scala 55:32]
  wire [1:0] _T_200; // @[LZD.scala 55:20]
  wire [2:0] _T_201; // @[Cat.scala 29:58]
  wire [2:0] _T_202; // @[convert.scala 21:22]
  wire [3:0] _T_203; // @[convert.scala 22:36]
  wire  _T_204; // @[Shift.scala 16:24]
  wire [1:0] _T_205; // @[Shift.scala 17:37]
  wire  _T_206; // @[Shift.scala 12:21]
  wire [1:0] _T_207; // @[Shift.scala 64:52]
  wire [3:0] _T_209; // @[Cat.scala 29:58]
  wire [3:0] _T_210; // @[Shift.scala 64:27]
  wire  _T_211; // @[Shift.scala 66:70]
  wire [2:0] _T_213; // @[Shift.scala 64:52]
  wire [3:0] _T_214; // @[Cat.scala 29:58]
  wire  _T_219; // @[convert.scala 25:26]
  wire [2:0] _T_221; // @[convert.scala 25:42]
  wire [3:0] _T_222; // @[Cat.scala 29:58]
  wire [5:0] _T_224; // @[convert.scala 29:56]
  wire  _T_225; // @[convert.scala 29:60]
  wire  _T_226; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_229; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [3:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_237; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_238; // @[PositFMA.scala 59:34]
  wire  _T_239; // @[PositFMA.scala 59:47]
  wire  _T_240; // @[PositFMA.scala 59:45]
  wire [5:0] _T_242; // @[Cat.scala 29:58]
  wire [5:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_243; // @[PositFMA.scala 60:34]
  wire  _T_244; // @[PositFMA.scala 60:47]
  wire  _T_245; // @[PositFMA.scala 60:45]
  wire [5:0] _T_247; // @[Cat.scala 29:58]
  wire [5:0] sigB; // @[PositFMA.scala 60:76]
  wire [11:0] _T_248; // @[PositFMA.scala 62:25]
  wire [11:0] sigP; // @[PositFMA.scala 62:33]
  wire [1:0] head2; // @[PositFMA.scala 63:28]
  wire  _T_249; // @[PositFMA.scala 64:31]
  wire  _T_250; // @[PositFMA.scala 64:25]
  wire  _T_251; // @[PositFMA.scala 64:42]
  wire  addTwo; // @[PositFMA.scala 64:35]
  wire  _T_252; // @[PositFMA.scala 66:23]
  wire  _T_253; // @[PositFMA.scala 66:49]
  wire  addOne; // @[PositFMA.scala 66:43]
  wire [1:0] _T_254; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 67:39]
  wire  mulSign; // @[PositFMA.scala 68:28]
  wire [4:0] _T_255; // @[PositFMA.scala 70:30]
  wire [4:0] _GEN_12; // @[PositFMA.scala 70:44]
  wire [4:0] _T_257; // @[PositFMA.scala 70:44]
  wire [4:0] mulScale; // @[PositFMA.scala 70:44]
  wire [9:0] _T_258; // @[PositFMA.scala 73:29]
  wire [8:0] _T_259; // @[PositFMA.scala 74:29]
  wire [9:0] _T_260; // @[PositFMA.scala 74:48]
  wire [9:0] mulSigTmp; // @[PositFMA.scala 71:22]
  wire  _T_262; // @[PositFMA.scala 78:39]
  wire  _T_263; // @[PositFMA.scala 78:43]
  wire [8:0] _T_264; // @[PositFMA.scala 79:39]
  wire [10:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [10:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [3:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [4:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [3:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_290; // @[PositFMA.scala 108:29]
  wire  _T_291; // @[PositFMA.scala 108:47]
  wire  _T_292; // @[PositFMA.scala 108:45]
  wire [10:0] extAddSig; // @[Cat.scala 29:58]
  wire [4:0] _GEN_13; // @[PositFMA.scala 112:39]
  wire  mulGreater; // @[PositFMA.scala 112:39]
  wire [4:0] greaterScale; // @[PositFMA.scala 113:26]
  wire [4:0] smallerScale; // @[PositFMA.scala 114:26]
  wire [4:0] _T_296; // @[PositFMA.scala 115:36]
  wire [4:0] scaleDiff; // @[PositFMA.scala 115:36]
  wire [10:0] greaterSig; // @[PositFMA.scala 116:26]
  wire [10:0] smallerSigTmp; // @[PositFMA.scala 117:26]
  wire [4:0] _T_297; // @[PositFMA.scala 118:69]
  wire  _T_298; // @[Shift.scala 39:24]
  wire [3:0] _T_299; // @[Shift.scala 40:44]
  wire [2:0] _T_300; // @[Shift.scala 90:30]
  wire [7:0] _T_301; // @[Shift.scala 90:48]
  wire  _T_302; // @[Shift.scala 90:57]
  wire [2:0] _GEN_14; // @[Shift.scala 90:39]
  wire [2:0] _T_303; // @[Shift.scala 90:39]
  wire  _T_304; // @[Shift.scala 12:21]
  wire  _T_305; // @[Shift.scala 12:21]
  wire [7:0] _T_307; // @[Bitwise.scala 71:12]
  wire [10:0] _T_308; // @[Cat.scala 29:58]
  wire [10:0] _T_309; // @[Shift.scala 91:22]
  wire [2:0] _T_310; // @[Shift.scala 92:77]
  wire [6:0] _T_311; // @[Shift.scala 90:30]
  wire [3:0] _T_312; // @[Shift.scala 90:48]
  wire  _T_313; // @[Shift.scala 90:57]
  wire [6:0] _GEN_15; // @[Shift.scala 90:39]
  wire [6:0] _T_314; // @[Shift.scala 90:39]
  wire  _T_315; // @[Shift.scala 12:21]
  wire  _T_316; // @[Shift.scala 12:21]
  wire [3:0] _T_318; // @[Bitwise.scala 71:12]
  wire [10:0] _T_319; // @[Cat.scala 29:58]
  wire [10:0] _T_320; // @[Shift.scala 91:22]
  wire [1:0] _T_321; // @[Shift.scala 92:77]
  wire [8:0] _T_322; // @[Shift.scala 90:30]
  wire [1:0] _T_323; // @[Shift.scala 90:48]
  wire  _T_324; // @[Shift.scala 90:57]
  wire [8:0] _GEN_16; // @[Shift.scala 90:39]
  wire [8:0] _T_325; // @[Shift.scala 90:39]
  wire  _T_326; // @[Shift.scala 12:21]
  wire  _T_327; // @[Shift.scala 12:21]
  wire [1:0] _T_329; // @[Bitwise.scala 71:12]
  wire [10:0] _T_330; // @[Cat.scala 29:58]
  wire [10:0] _T_331; // @[Shift.scala 91:22]
  wire  _T_332; // @[Shift.scala 92:77]
  wire [9:0] _T_333; // @[Shift.scala 90:30]
  wire  _T_334; // @[Shift.scala 90:48]
  wire [9:0] _GEN_17; // @[Shift.scala 90:39]
  wire [9:0] _T_336; // @[Shift.scala 90:39]
  wire  _T_338; // @[Shift.scala 12:21]
  wire [10:0] _T_339; // @[Cat.scala 29:58]
  wire [10:0] _T_340; // @[Shift.scala 91:22]
  wire [10:0] _T_343; // @[Bitwise.scala 71:12]
  wire [10:0] smallerSig; // @[Shift.scala 39:10]
  wire [11:0] rawSumSig; // @[PositFMA.scala 119:34]
  wire  _T_344; // @[PositFMA.scala 120:42]
  wire  _T_345; // @[PositFMA.scala 120:46]
  wire  _T_346; // @[PositFMA.scala 120:79]
  wire  sumSign; // @[PositFMA.scala 120:63]
  wire [10:0] _T_348; // @[PositFMA.scala 121:50]
  wire [11:0] signSumSig; // @[Cat.scala 29:58]
  wire [10:0] _T_349; // @[PositFMA.scala 126:33]
  wire [10:0] _T_350; // @[PositFMA.scala 126:68]
  wire [10:0] sumXor; // @[PositFMA.scala 126:51]
  wire [7:0] _T_351; // @[LZD.scala 43:32]
  wire [3:0] _T_352; // @[LZD.scala 43:32]
  wire [1:0] _T_353; // @[LZD.scala 43:32]
  wire  _T_354; // @[LZD.scala 39:14]
  wire  _T_355; // @[LZD.scala 39:21]
  wire  _T_356; // @[LZD.scala 39:30]
  wire  _T_357; // @[LZD.scala 39:27]
  wire  _T_358; // @[LZD.scala 39:25]
  wire [1:0] _T_359; // @[Cat.scala 29:58]
  wire [1:0] _T_360; // @[LZD.scala 44:32]
  wire  _T_361; // @[LZD.scala 39:14]
  wire  _T_362; // @[LZD.scala 39:21]
  wire  _T_363; // @[LZD.scala 39:30]
  wire  _T_364; // @[LZD.scala 39:27]
  wire  _T_365; // @[LZD.scala 39:25]
  wire [1:0] _T_366; // @[Cat.scala 29:58]
  wire  _T_367; // @[Shift.scala 12:21]
  wire  _T_368; // @[Shift.scala 12:21]
  wire  _T_369; // @[LZD.scala 49:16]
  wire  _T_370; // @[LZD.scala 49:27]
  wire  _T_371; // @[LZD.scala 49:25]
  wire  _T_372; // @[LZD.scala 49:47]
  wire  _T_373; // @[LZD.scala 49:59]
  wire  _T_374; // @[LZD.scala 49:35]
  wire [2:0] _T_376; // @[Cat.scala 29:58]
  wire [3:0] _T_377; // @[LZD.scala 44:32]
  wire [1:0] _T_378; // @[LZD.scala 43:32]
  wire  _T_379; // @[LZD.scala 39:14]
  wire  _T_380; // @[LZD.scala 39:21]
  wire  _T_381; // @[LZD.scala 39:30]
  wire  _T_382; // @[LZD.scala 39:27]
  wire  _T_383; // @[LZD.scala 39:25]
  wire [1:0] _T_384; // @[Cat.scala 29:58]
  wire [1:0] _T_385; // @[LZD.scala 44:32]
  wire  _T_386; // @[LZD.scala 39:14]
  wire  _T_387; // @[LZD.scala 39:21]
  wire  _T_388; // @[LZD.scala 39:30]
  wire  _T_389; // @[LZD.scala 39:27]
  wire  _T_390; // @[LZD.scala 39:25]
  wire [1:0] _T_391; // @[Cat.scala 29:58]
  wire  _T_392; // @[Shift.scala 12:21]
  wire  _T_393; // @[Shift.scala 12:21]
  wire  _T_394; // @[LZD.scala 49:16]
  wire  _T_395; // @[LZD.scala 49:27]
  wire  _T_396; // @[LZD.scala 49:25]
  wire  _T_397; // @[LZD.scala 49:47]
  wire  _T_398; // @[LZD.scala 49:59]
  wire  _T_399; // @[LZD.scala 49:35]
  wire [2:0] _T_401; // @[Cat.scala 29:58]
  wire  _T_402; // @[Shift.scala 12:21]
  wire  _T_403; // @[Shift.scala 12:21]
  wire  _T_404; // @[LZD.scala 49:16]
  wire  _T_405; // @[LZD.scala 49:27]
  wire  _T_406; // @[LZD.scala 49:25]
  wire [1:0] _T_407; // @[LZD.scala 49:47]
  wire [1:0] _T_408; // @[LZD.scala 49:59]
  wire [1:0] _T_409; // @[LZD.scala 49:35]
  wire [3:0] _T_411; // @[Cat.scala 29:58]
  wire [2:0] _T_412; // @[LZD.scala 44:32]
  wire [1:0] _T_413; // @[LZD.scala 43:32]
  wire  _T_414; // @[LZD.scala 39:14]
  wire  _T_415; // @[LZD.scala 39:21]
  wire  _T_416; // @[LZD.scala 39:30]
  wire  _T_417; // @[LZD.scala 39:27]
  wire  _T_418; // @[LZD.scala 39:25]
  wire [1:0] _T_419; // @[Cat.scala 29:58]
  wire  _T_420; // @[LZD.scala 44:32]
  wire  _T_422; // @[Shift.scala 12:21]
  wire  _T_424; // @[LZD.scala 55:32]
  wire  _T_425; // @[LZD.scala 55:20]
  wire  _T_427; // @[Shift.scala 12:21]
  wire [2:0] _T_429; // @[Cat.scala 29:58]
  wire [2:0] _T_430; // @[LZD.scala 55:32]
  wire [2:0] _T_431; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [3:0] shiftValue; // @[PositFMA.scala 128:24]
  wire [9:0] _T_432; // @[PositFMA.scala 129:38]
  wire  _T_433; // @[Shift.scala 16:24]
  wire  _T_435; // @[Shift.scala 12:21]
  wire [1:0] _T_436; // @[Shift.scala 64:52]
  wire [9:0] _T_438; // @[Cat.scala 29:58]
  wire [9:0] _T_439; // @[Shift.scala 64:27]
  wire [2:0] _T_440; // @[Shift.scala 66:70]
  wire  _T_441; // @[Shift.scala 12:21]
  wire [5:0] _T_442; // @[Shift.scala 64:52]
  wire [9:0] _T_444; // @[Cat.scala 29:58]
  wire [9:0] _T_445; // @[Shift.scala 64:27]
  wire [1:0] _T_446; // @[Shift.scala 66:70]
  wire  _T_447; // @[Shift.scala 12:21]
  wire [7:0] _T_448; // @[Shift.scala 64:52]
  wire [9:0] _T_450; // @[Cat.scala 29:58]
  wire [9:0] _T_451; // @[Shift.scala 64:27]
  wire  _T_452; // @[Shift.scala 66:70]
  wire [8:0] _T_454; // @[Shift.scala 64:52]
  wire [9:0] _T_455; // @[Cat.scala 29:58]
  wire [9:0] _T_456; // @[Shift.scala 64:27]
  wire [9:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [4:0] _T_458; // @[PositFMA.scala 132:36]
  wire [4:0] _T_459; // @[PositFMA.scala 132:36]
  wire [4:0] _T_460; // @[Cat.scala 29:58]
  wire [4:0] _T_461; // @[PositFMA.scala 132:61]
  wire [4:0] _T_463; // @[PositFMA.scala 132:42]
  wire [4:0] sumScale; // @[PositFMA.scala 132:42]
  wire [3:0] sumFrac; // @[PositFMA.scala 133:41]
  wire [5:0] grsTmp; // @[PositFMA.scala 136:41]
  wire [1:0] _T_464; // @[PositFMA.scala 139:40]
  wire [3:0] _T_465; // @[PositFMA.scala 139:56]
  wire  _T_466; // @[PositFMA.scala 139:60]
  wire  underflow; // @[PositFMA.scala 146:32]
  wire  overflow; // @[PositFMA.scala 147:32]
  wire  _T_467; // @[PositFMA.scala 156:32]
  wire  decF_isZero; // @[PositFMA.scala 156:20]
  wire [4:0] _T_469; // @[Mux.scala 87:16]
  wire [4:0] _T_470; // @[Mux.scala 87:16]
  wire [3:0] _GEN_18; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  wire [3:0] decF_scale; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  wire  _T_472; // @[convert.scala 49:36]
  wire [3:0] _T_474; // @[convert.scala 50:36]
  wire [3:0] _T_475; // @[convert.scala 50:36]
  wire [3:0] _T_476; // @[convert.scala 50:28]
  wire  _T_477; // @[convert.scala 51:31]
  wire  _T_478; // @[convert.scala 53:34]
  wire [8:0] _T_481; // @[Cat.scala 29:58]
  wire [3:0] _T_482; // @[Shift.scala 39:17]
  wire  _T_483; // @[Shift.scala 39:24]
  wire  _T_485; // @[Shift.scala 90:30]
  wire [7:0] _T_486; // @[Shift.scala 90:48]
  wire  _T_487; // @[Shift.scala 90:57]
  wire  _T_488; // @[Shift.scala 90:39]
  wire  _T_489; // @[Shift.scala 12:21]
  wire  _T_490; // @[Shift.scala 12:21]
  wire [7:0] _T_492; // @[Bitwise.scala 71:12]
  wire [8:0] _T_493; // @[Cat.scala 29:58]
  wire [8:0] _T_494; // @[Shift.scala 91:22]
  wire [2:0] _T_495; // @[Shift.scala 92:77]
  wire [4:0] _T_496; // @[Shift.scala 90:30]
  wire [3:0] _T_497; // @[Shift.scala 90:48]
  wire  _T_498; // @[Shift.scala 90:57]
  wire [4:0] _GEN_19; // @[Shift.scala 90:39]
  wire [4:0] _T_499; // @[Shift.scala 90:39]
  wire  _T_500; // @[Shift.scala 12:21]
  wire  _T_501; // @[Shift.scala 12:21]
  wire [3:0] _T_503; // @[Bitwise.scala 71:12]
  wire [8:0] _T_504; // @[Cat.scala 29:58]
  wire [8:0] _T_505; // @[Shift.scala 91:22]
  wire [1:0] _T_506; // @[Shift.scala 92:77]
  wire [6:0] _T_507; // @[Shift.scala 90:30]
  wire [1:0] _T_508; // @[Shift.scala 90:48]
  wire  _T_509; // @[Shift.scala 90:57]
  wire [6:0] _GEN_20; // @[Shift.scala 90:39]
  wire [6:0] _T_510; // @[Shift.scala 90:39]
  wire  _T_511; // @[Shift.scala 12:21]
  wire  _T_512; // @[Shift.scala 12:21]
  wire [1:0] _T_514; // @[Bitwise.scala 71:12]
  wire [8:0] _T_515; // @[Cat.scala 29:58]
  wire [8:0] _T_516; // @[Shift.scala 91:22]
  wire  _T_517; // @[Shift.scala 92:77]
  wire [7:0] _T_518; // @[Shift.scala 90:30]
  wire  _T_519; // @[Shift.scala 90:48]
  wire [7:0] _GEN_21; // @[Shift.scala 90:39]
  wire [7:0] _T_521; // @[Shift.scala 90:39]
  wire  _T_523; // @[Shift.scala 12:21]
  wire [8:0] _T_524; // @[Cat.scala 29:58]
  wire [8:0] _T_525; // @[Shift.scala 91:22]
  wire [8:0] _T_528; // @[Bitwise.scala 71:12]
  wire [8:0] _T_529; // @[Shift.scala 39:10]
  wire  _T_530; // @[convert.scala 55:31]
  wire  _T_531; // @[convert.scala 56:31]
  wire  _T_532; // @[convert.scala 57:31]
  wire  _T_533; // @[convert.scala 58:31]
  wire [5:0] _T_534; // @[convert.scala 59:69]
  wire  _T_535; // @[convert.scala 59:81]
  wire  _T_536; // @[convert.scala 59:50]
  wire  _T_538; // @[convert.scala 60:81]
  wire  _T_539; // @[convert.scala 61:44]
  wire  _T_540; // @[convert.scala 61:52]
  wire  _T_541; // @[convert.scala 61:36]
  wire  _T_542; // @[convert.scala 62:63]
  wire  _T_543; // @[convert.scala 62:103]
  wire  _T_544; // @[convert.scala 62:60]
  wire [5:0] _GEN_22; // @[convert.scala 63:56]
  wire [5:0] _T_547; // @[convert.scala 63:56]
  wire [6:0] _T_548; // @[Cat.scala 29:58]
  reg  _T_552; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [6:0] _T_556; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{6'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{6'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[6]; // @[convert.scala 18:24]
  assign _T_14 = realA[5]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[5:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[4:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[4:1]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[3:2]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20 != 2'h0; // @[LZD.scala 39:14]
  assign _T_22 = _T_20[1]; // @[LZD.scala 39:21]
  assign _T_23 = _T_20[0]; // @[LZD.scala 39:30]
  assign _T_24 = ~ _T_23; // @[LZD.scala 39:27]
  assign _T_25 = _T_22 | _T_24; // @[LZD.scala 39:25]
  assign _T_26 = {_T_21,_T_25}; // @[Cat.scala 29:58]
  assign _T_27 = _T_19[1:0]; // @[LZD.scala 44:32]
  assign _T_28 = _T_27 != 2'h0; // @[LZD.scala 39:14]
  assign _T_29 = _T_27[1]; // @[LZD.scala 39:21]
  assign _T_30 = _T_27[0]; // @[LZD.scala 39:30]
  assign _T_31 = ~ _T_30; // @[LZD.scala 39:27]
  assign _T_32 = _T_29 | _T_31; // @[LZD.scala 39:25]
  assign _T_33 = {_T_28,_T_32}; // @[Cat.scala 29:58]
  assign _T_34 = _T_26[1]; // @[Shift.scala 12:21]
  assign _T_35 = _T_33[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_34 | _T_35; // @[LZD.scala 49:16]
  assign _T_37 = ~ _T_35; // @[LZD.scala 49:27]
  assign _T_38 = _T_34 | _T_37; // @[LZD.scala 49:25]
  assign _T_39 = _T_26[0:0]; // @[LZD.scala 49:47]
  assign _T_40 = _T_33[0:0]; // @[LZD.scala 49:59]
  assign _T_41 = _T_34 ? _T_39 : _T_40; // @[LZD.scala 49:35]
  assign _T_43 = {_T_36,_T_38,_T_41}; // @[Cat.scala 29:58]
  assign _T_44 = _T_18[0:0]; // @[LZD.scala 44:32]
  assign _T_46 = _T_43[2]; // @[Shift.scala 12:21]
  assign _T_48 = {1'h1,_T_44}; // @[Cat.scala 29:58]
  assign _T_49 = _T_43[1:0]; // @[LZD.scala 55:32]
  assign _T_50 = _T_46 ? _T_49 : _T_48; // @[LZD.scala 55:20]
  assign _T_51 = {_T_46,_T_50}; // @[Cat.scala 29:58]
  assign _T_52 = ~ _T_51; // @[convert.scala 21:22]
  assign _T_53 = realA[3:0]; // @[convert.scala 22:36]
  assign _T_54 = _T_52 < 3'h4; // @[Shift.scala 16:24]
  assign _T_55 = _T_52[1:0]; // @[Shift.scala 17:37]
  assign _T_56 = _T_55[1]; // @[Shift.scala 12:21]
  assign _T_57 = _T_53[1:0]; // @[Shift.scala 64:52]
  assign _T_59 = {_T_57,2'h0}; // @[Cat.scala 29:58]
  assign _T_60 = _T_56 ? _T_59 : _T_53; // @[Shift.scala 64:27]
  assign _T_61 = _T_55[0:0]; // @[Shift.scala 66:70]
  assign _T_63 = _T_60[2:0]; // @[Shift.scala 64:52]
  assign _T_64 = {_T_63,1'h0}; // @[Cat.scala 29:58]
  assign _T_65 = _T_61 ? _T_64 : _T_60; // @[Shift.scala 64:27]
  assign decA_fraction = _T_54 ? _T_65 : 4'h0; // @[Shift.scala 16:10]
  assign _T_69 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_71 = _T_15 ? _T_52 : _T_51; // @[convert.scala 25:42]
  assign _T_72 = {_T_69,_T_71}; // @[Cat.scala 29:58]
  assign _T_74 = realA[5:0]; // @[convert.scala 29:56]
  assign _T_75 = _T_74 != 6'h0; // @[convert.scala 29:60]
  assign _T_76 = ~ _T_75; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_76; // @[convert.scala 29:39]
  assign _T_79 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_79 & _T_76; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_72); // @[convert.scala 32:24]
  assign _T_88 = io_B[6]; // @[convert.scala 18:24]
  assign _T_89 = io_B[5]; // @[convert.scala 18:40]
  assign _T_90 = _T_88 ^ _T_89; // @[convert.scala 18:36]
  assign _T_91 = io_B[5:1]; // @[convert.scala 19:24]
  assign _T_92 = io_B[4:0]; // @[convert.scala 19:43]
  assign _T_93 = _T_91 ^ _T_92; // @[convert.scala 19:39]
  assign _T_94 = _T_93[4:1]; // @[LZD.scala 43:32]
  assign _T_95 = _T_94[3:2]; // @[LZD.scala 43:32]
  assign _T_96 = _T_95 != 2'h0; // @[LZD.scala 39:14]
  assign _T_97 = _T_95[1]; // @[LZD.scala 39:21]
  assign _T_98 = _T_95[0]; // @[LZD.scala 39:30]
  assign _T_99 = ~ _T_98; // @[LZD.scala 39:27]
  assign _T_100 = _T_97 | _T_99; // @[LZD.scala 39:25]
  assign _T_101 = {_T_96,_T_100}; // @[Cat.scala 29:58]
  assign _T_102 = _T_94[1:0]; // @[LZD.scala 44:32]
  assign _T_103 = _T_102 != 2'h0; // @[LZD.scala 39:14]
  assign _T_104 = _T_102[1]; // @[LZD.scala 39:21]
  assign _T_105 = _T_102[0]; // @[LZD.scala 39:30]
  assign _T_106 = ~ _T_105; // @[LZD.scala 39:27]
  assign _T_107 = _T_104 | _T_106; // @[LZD.scala 39:25]
  assign _T_108 = {_T_103,_T_107}; // @[Cat.scala 29:58]
  assign _T_109 = _T_101[1]; // @[Shift.scala 12:21]
  assign _T_110 = _T_108[1]; // @[Shift.scala 12:21]
  assign _T_111 = _T_109 | _T_110; // @[LZD.scala 49:16]
  assign _T_112 = ~ _T_110; // @[LZD.scala 49:27]
  assign _T_113 = _T_109 | _T_112; // @[LZD.scala 49:25]
  assign _T_114 = _T_101[0:0]; // @[LZD.scala 49:47]
  assign _T_115 = _T_108[0:0]; // @[LZD.scala 49:59]
  assign _T_116 = _T_109 ? _T_114 : _T_115; // @[LZD.scala 49:35]
  assign _T_118 = {_T_111,_T_113,_T_116}; // @[Cat.scala 29:58]
  assign _T_119 = _T_93[0:0]; // @[LZD.scala 44:32]
  assign _T_121 = _T_118[2]; // @[Shift.scala 12:21]
  assign _T_123 = {1'h1,_T_119}; // @[Cat.scala 29:58]
  assign _T_124 = _T_118[1:0]; // @[LZD.scala 55:32]
  assign _T_125 = _T_121 ? _T_124 : _T_123; // @[LZD.scala 55:20]
  assign _T_126 = {_T_121,_T_125}; // @[Cat.scala 29:58]
  assign _T_127 = ~ _T_126; // @[convert.scala 21:22]
  assign _T_128 = io_B[3:0]; // @[convert.scala 22:36]
  assign _T_129 = _T_127 < 3'h4; // @[Shift.scala 16:24]
  assign _T_130 = _T_127[1:0]; // @[Shift.scala 17:37]
  assign _T_131 = _T_130[1]; // @[Shift.scala 12:21]
  assign _T_132 = _T_128[1:0]; // @[Shift.scala 64:52]
  assign _T_134 = {_T_132,2'h0}; // @[Cat.scala 29:58]
  assign _T_135 = _T_131 ? _T_134 : _T_128; // @[Shift.scala 64:27]
  assign _T_136 = _T_130[0:0]; // @[Shift.scala 66:70]
  assign _T_138 = _T_135[2:0]; // @[Shift.scala 64:52]
  assign _T_139 = {_T_138,1'h0}; // @[Cat.scala 29:58]
  assign _T_140 = _T_136 ? _T_139 : _T_135; // @[Shift.scala 64:27]
  assign decB_fraction = _T_129 ? _T_140 : 4'h0; // @[Shift.scala 16:10]
  assign _T_144 = _T_90 == 1'h0; // @[convert.scala 25:26]
  assign _T_146 = _T_90 ? _T_127 : _T_126; // @[convert.scala 25:42]
  assign _T_147 = {_T_144,_T_146}; // @[Cat.scala 29:58]
  assign _T_149 = io_B[5:0]; // @[convert.scala 29:56]
  assign _T_150 = _T_149 != 6'h0; // @[convert.scala 29:60]
  assign _T_151 = ~ _T_150; // @[convert.scala 29:41]
  assign decB_isNaR = _T_88 & _T_151; // @[convert.scala 29:39]
  assign _T_154 = _T_88 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_154 & _T_151; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_147); // @[convert.scala 32:24]
  assign _T_163 = realC[6]; // @[convert.scala 18:24]
  assign _T_164 = realC[5]; // @[convert.scala 18:40]
  assign _T_165 = _T_163 ^ _T_164; // @[convert.scala 18:36]
  assign _T_166 = realC[5:1]; // @[convert.scala 19:24]
  assign _T_167 = realC[4:0]; // @[convert.scala 19:43]
  assign _T_168 = _T_166 ^ _T_167; // @[convert.scala 19:39]
  assign _T_169 = _T_168[4:1]; // @[LZD.scala 43:32]
  assign _T_170 = _T_169[3:2]; // @[LZD.scala 43:32]
  assign _T_171 = _T_170 != 2'h0; // @[LZD.scala 39:14]
  assign _T_172 = _T_170[1]; // @[LZD.scala 39:21]
  assign _T_173 = _T_170[0]; // @[LZD.scala 39:30]
  assign _T_174 = ~ _T_173; // @[LZD.scala 39:27]
  assign _T_175 = _T_172 | _T_174; // @[LZD.scala 39:25]
  assign _T_176 = {_T_171,_T_175}; // @[Cat.scala 29:58]
  assign _T_177 = _T_169[1:0]; // @[LZD.scala 44:32]
  assign _T_178 = _T_177 != 2'h0; // @[LZD.scala 39:14]
  assign _T_179 = _T_177[1]; // @[LZD.scala 39:21]
  assign _T_180 = _T_177[0]; // @[LZD.scala 39:30]
  assign _T_181 = ~ _T_180; // @[LZD.scala 39:27]
  assign _T_182 = _T_179 | _T_181; // @[LZD.scala 39:25]
  assign _T_183 = {_T_178,_T_182}; // @[Cat.scala 29:58]
  assign _T_184 = _T_176[1]; // @[Shift.scala 12:21]
  assign _T_185 = _T_183[1]; // @[Shift.scala 12:21]
  assign _T_186 = _T_184 | _T_185; // @[LZD.scala 49:16]
  assign _T_187 = ~ _T_185; // @[LZD.scala 49:27]
  assign _T_188 = _T_184 | _T_187; // @[LZD.scala 49:25]
  assign _T_189 = _T_176[0:0]; // @[LZD.scala 49:47]
  assign _T_190 = _T_183[0:0]; // @[LZD.scala 49:59]
  assign _T_191 = _T_184 ? _T_189 : _T_190; // @[LZD.scala 49:35]
  assign _T_193 = {_T_186,_T_188,_T_191}; // @[Cat.scala 29:58]
  assign _T_194 = _T_168[0:0]; // @[LZD.scala 44:32]
  assign _T_196 = _T_193[2]; // @[Shift.scala 12:21]
  assign _T_198 = {1'h1,_T_194}; // @[Cat.scala 29:58]
  assign _T_199 = _T_193[1:0]; // @[LZD.scala 55:32]
  assign _T_200 = _T_196 ? _T_199 : _T_198; // @[LZD.scala 55:20]
  assign _T_201 = {_T_196,_T_200}; // @[Cat.scala 29:58]
  assign _T_202 = ~ _T_201; // @[convert.scala 21:22]
  assign _T_203 = realC[3:0]; // @[convert.scala 22:36]
  assign _T_204 = _T_202 < 3'h4; // @[Shift.scala 16:24]
  assign _T_205 = _T_202[1:0]; // @[Shift.scala 17:37]
  assign _T_206 = _T_205[1]; // @[Shift.scala 12:21]
  assign _T_207 = _T_203[1:0]; // @[Shift.scala 64:52]
  assign _T_209 = {_T_207,2'h0}; // @[Cat.scala 29:58]
  assign _T_210 = _T_206 ? _T_209 : _T_203; // @[Shift.scala 64:27]
  assign _T_211 = _T_205[0:0]; // @[Shift.scala 66:70]
  assign _T_213 = _T_210[2:0]; // @[Shift.scala 64:52]
  assign _T_214 = {_T_213,1'h0}; // @[Cat.scala 29:58]
  assign _T_219 = _T_165 == 1'h0; // @[convert.scala 25:26]
  assign _T_221 = _T_165 ? _T_202 : _T_201; // @[convert.scala 25:42]
  assign _T_222 = {_T_219,_T_221}; // @[Cat.scala 29:58]
  assign _T_224 = realC[5:0]; // @[convert.scala 29:56]
  assign _T_225 = _T_224 != 6'h0; // @[convert.scala 29:60]
  assign _T_226 = ~ _T_225; // @[convert.scala 29:41]
  assign decC_isNaR = _T_163 & _T_226; // @[convert.scala 29:39]
  assign _T_229 = _T_163 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_229 & _T_226; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_222); // @[convert.scala 32:24]
  assign _T_237 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_237 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_238 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_239 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_240 = _T_238 & _T_239; // @[PositFMA.scala 59:45]
  assign _T_242 = {_T_13,_T_240,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_242); // @[PositFMA.scala 59:76]
  assign _T_243 = ~ _T_88; // @[PositFMA.scala 60:34]
  assign _T_244 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_245 = _T_243 & _T_244; // @[PositFMA.scala 60:45]
  assign _T_247 = {_T_88,_T_245,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_247); // @[PositFMA.scala 60:76]
  assign _T_248 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 62:25]
  assign sigP = $unsigned(_T_248); // @[PositFMA.scala 62:33]
  assign head2 = sigP[11:10]; // @[PositFMA.scala 63:28]
  assign _T_249 = head2[1]; // @[PositFMA.scala 64:31]
  assign _T_250 = ~ _T_249; // @[PositFMA.scala 64:25]
  assign _T_251 = head2[0]; // @[PositFMA.scala 64:42]
  assign addTwo = _T_250 & _T_251; // @[PositFMA.scala 64:35]
  assign _T_252 = sigP[11]; // @[PositFMA.scala 66:23]
  assign _T_253 = sigP[9]; // @[PositFMA.scala 66:49]
  assign addOne = _T_252 ^ _T_253; // @[PositFMA.scala 66:43]
  assign _T_254 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_254)}; // @[PositFMA.scala 67:39]
  assign mulSign = sigP[11:11]; // @[PositFMA.scala 68:28]
  assign _T_255 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 70:30]
  assign _GEN_12 = {{2{expBias[2]}},expBias}; // @[PositFMA.scala 70:44]
  assign _T_257 = $signed(_T_255) + $signed(_GEN_12); // @[PositFMA.scala 70:44]
  assign mulScale = $signed(_T_257); // @[PositFMA.scala 70:44]
  assign _T_258 = sigP[9:0]; // @[PositFMA.scala 73:29]
  assign _T_259 = sigP[8:0]; // @[PositFMA.scala 74:29]
  assign _T_260 = {_T_259, 1'h0}; // @[PositFMA.scala 74:48]
  assign mulSigTmp = addOne ? _T_258 : _T_260; // @[PositFMA.scala 71:22]
  assign _T_262 = mulSigTmp[9:9]; // @[PositFMA.scala 78:39]
  assign _T_263 = _T_262 | addTwo; // @[PositFMA.scala 78:43]
  assign _T_264 = mulSigTmp[8:0]; // @[PositFMA.scala 79:39]
  assign mulSig = {mulSign,_T_263,_T_264}; // @[Cat.scala 29:58]
  assign _T_290 = ~ addSign_phase2; // @[PositFMA.scala 108:29]
  assign _T_291 = ~ addZero_phase2; // @[PositFMA.scala 108:47]
  assign _T_292 = _T_290 & _T_291; // @[PositFMA.scala 108:45]
  assign extAddSig = {addSign_phase2,_T_292,addFrac_phase2,5'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[3]}},addScale_phase2}; // @[PositFMA.scala 112:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 112:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[3]}},addScale_phase2}); // @[PositFMA.scala 113:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[3]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 114:26]
  assign _T_296 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 115:36]
  assign scaleDiff = $signed(_T_296); // @[PositFMA.scala 115:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 116:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 117:26]
  assign _T_297 = $unsigned(scaleDiff); // @[PositFMA.scala 118:69]
  assign _T_298 = _T_297 < 5'hb; // @[Shift.scala 39:24]
  assign _T_299 = _T_297[3:0]; // @[Shift.scala 40:44]
  assign _T_300 = smallerSigTmp[10:8]; // @[Shift.scala 90:30]
  assign _T_301 = smallerSigTmp[7:0]; // @[Shift.scala 90:48]
  assign _T_302 = _T_301 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{2'd0}, _T_302}; // @[Shift.scala 90:39]
  assign _T_303 = _T_300 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_304 = _T_299[3]; // @[Shift.scala 12:21]
  assign _T_305 = smallerSigTmp[10]; // @[Shift.scala 12:21]
  assign _T_307 = _T_305 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_308 = {_T_307,_T_303}; // @[Cat.scala 29:58]
  assign _T_309 = _T_304 ? _T_308 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_310 = _T_299[2:0]; // @[Shift.scala 92:77]
  assign _T_311 = _T_309[10:4]; // @[Shift.scala 90:30]
  assign _T_312 = _T_309[3:0]; // @[Shift.scala 90:48]
  assign _T_313 = _T_312 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{6'd0}, _T_313}; // @[Shift.scala 90:39]
  assign _T_314 = _T_311 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_315 = _T_310[2]; // @[Shift.scala 12:21]
  assign _T_316 = _T_309[10]; // @[Shift.scala 12:21]
  assign _T_318 = _T_316 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_319 = {_T_318,_T_314}; // @[Cat.scala 29:58]
  assign _T_320 = _T_315 ? _T_319 : _T_309; // @[Shift.scala 91:22]
  assign _T_321 = _T_310[1:0]; // @[Shift.scala 92:77]
  assign _T_322 = _T_320[10:2]; // @[Shift.scala 90:30]
  assign _T_323 = _T_320[1:0]; // @[Shift.scala 90:48]
  assign _T_324 = _T_323 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_16 = {{8'd0}, _T_324}; // @[Shift.scala 90:39]
  assign _T_325 = _T_322 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_326 = _T_321[1]; // @[Shift.scala 12:21]
  assign _T_327 = _T_320[10]; // @[Shift.scala 12:21]
  assign _T_329 = _T_327 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_330 = {_T_329,_T_325}; // @[Cat.scala 29:58]
  assign _T_331 = _T_326 ? _T_330 : _T_320; // @[Shift.scala 91:22]
  assign _T_332 = _T_321[0:0]; // @[Shift.scala 92:77]
  assign _T_333 = _T_331[10:1]; // @[Shift.scala 90:30]
  assign _T_334 = _T_331[0:0]; // @[Shift.scala 90:48]
  assign _GEN_17 = {{9'd0}, _T_334}; // @[Shift.scala 90:39]
  assign _T_336 = _T_333 | _GEN_17; // @[Shift.scala 90:39]
  assign _T_338 = _T_331[10]; // @[Shift.scala 12:21]
  assign _T_339 = {_T_338,_T_336}; // @[Cat.scala 29:58]
  assign _T_340 = _T_332 ? _T_339 : _T_331; // @[Shift.scala 91:22]
  assign _T_343 = _T_305 ? 11'h7ff : 11'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_298 ? _T_340 : _T_343; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 119:34]
  assign _T_344 = mulSig_phase2[10:10]; // @[PositFMA.scala 120:42]
  assign _T_345 = _T_344 ^ addSign_phase2; // @[PositFMA.scala 120:46]
  assign _T_346 = rawSumSig[11:11]; // @[PositFMA.scala 120:79]
  assign sumSign = _T_345 ^ _T_346; // @[PositFMA.scala 120:63]
  assign _T_348 = greaterSig + smallerSig; // @[PositFMA.scala 121:50]
  assign signSumSig = {sumSign,_T_348}; // @[Cat.scala 29:58]
  assign _T_349 = signSumSig[11:1]; // @[PositFMA.scala 126:33]
  assign _T_350 = signSumSig[10:0]; // @[PositFMA.scala 126:68]
  assign sumXor = _T_349 ^ _T_350; // @[PositFMA.scala 126:51]
  assign _T_351 = sumXor[10:3]; // @[LZD.scala 43:32]
  assign _T_352 = _T_351[7:4]; // @[LZD.scala 43:32]
  assign _T_353 = _T_352[3:2]; // @[LZD.scala 43:32]
  assign _T_354 = _T_353 != 2'h0; // @[LZD.scala 39:14]
  assign _T_355 = _T_353[1]; // @[LZD.scala 39:21]
  assign _T_356 = _T_353[0]; // @[LZD.scala 39:30]
  assign _T_357 = ~ _T_356; // @[LZD.scala 39:27]
  assign _T_358 = _T_355 | _T_357; // @[LZD.scala 39:25]
  assign _T_359 = {_T_354,_T_358}; // @[Cat.scala 29:58]
  assign _T_360 = _T_352[1:0]; // @[LZD.scala 44:32]
  assign _T_361 = _T_360 != 2'h0; // @[LZD.scala 39:14]
  assign _T_362 = _T_360[1]; // @[LZD.scala 39:21]
  assign _T_363 = _T_360[0]; // @[LZD.scala 39:30]
  assign _T_364 = ~ _T_363; // @[LZD.scala 39:27]
  assign _T_365 = _T_362 | _T_364; // @[LZD.scala 39:25]
  assign _T_366 = {_T_361,_T_365}; // @[Cat.scala 29:58]
  assign _T_367 = _T_359[1]; // @[Shift.scala 12:21]
  assign _T_368 = _T_366[1]; // @[Shift.scala 12:21]
  assign _T_369 = _T_367 | _T_368; // @[LZD.scala 49:16]
  assign _T_370 = ~ _T_368; // @[LZD.scala 49:27]
  assign _T_371 = _T_367 | _T_370; // @[LZD.scala 49:25]
  assign _T_372 = _T_359[0:0]; // @[LZD.scala 49:47]
  assign _T_373 = _T_366[0:0]; // @[LZD.scala 49:59]
  assign _T_374 = _T_367 ? _T_372 : _T_373; // @[LZD.scala 49:35]
  assign _T_376 = {_T_369,_T_371,_T_374}; // @[Cat.scala 29:58]
  assign _T_377 = _T_351[3:0]; // @[LZD.scala 44:32]
  assign _T_378 = _T_377[3:2]; // @[LZD.scala 43:32]
  assign _T_379 = _T_378 != 2'h0; // @[LZD.scala 39:14]
  assign _T_380 = _T_378[1]; // @[LZD.scala 39:21]
  assign _T_381 = _T_378[0]; // @[LZD.scala 39:30]
  assign _T_382 = ~ _T_381; // @[LZD.scala 39:27]
  assign _T_383 = _T_380 | _T_382; // @[LZD.scala 39:25]
  assign _T_384 = {_T_379,_T_383}; // @[Cat.scala 29:58]
  assign _T_385 = _T_377[1:0]; // @[LZD.scala 44:32]
  assign _T_386 = _T_385 != 2'h0; // @[LZD.scala 39:14]
  assign _T_387 = _T_385[1]; // @[LZD.scala 39:21]
  assign _T_388 = _T_385[0]; // @[LZD.scala 39:30]
  assign _T_389 = ~ _T_388; // @[LZD.scala 39:27]
  assign _T_390 = _T_387 | _T_389; // @[LZD.scala 39:25]
  assign _T_391 = {_T_386,_T_390}; // @[Cat.scala 29:58]
  assign _T_392 = _T_384[1]; // @[Shift.scala 12:21]
  assign _T_393 = _T_391[1]; // @[Shift.scala 12:21]
  assign _T_394 = _T_392 | _T_393; // @[LZD.scala 49:16]
  assign _T_395 = ~ _T_393; // @[LZD.scala 49:27]
  assign _T_396 = _T_392 | _T_395; // @[LZD.scala 49:25]
  assign _T_397 = _T_384[0:0]; // @[LZD.scala 49:47]
  assign _T_398 = _T_391[0:0]; // @[LZD.scala 49:59]
  assign _T_399 = _T_392 ? _T_397 : _T_398; // @[LZD.scala 49:35]
  assign _T_401 = {_T_394,_T_396,_T_399}; // @[Cat.scala 29:58]
  assign _T_402 = _T_376[2]; // @[Shift.scala 12:21]
  assign _T_403 = _T_401[2]; // @[Shift.scala 12:21]
  assign _T_404 = _T_402 | _T_403; // @[LZD.scala 49:16]
  assign _T_405 = ~ _T_403; // @[LZD.scala 49:27]
  assign _T_406 = _T_402 | _T_405; // @[LZD.scala 49:25]
  assign _T_407 = _T_376[1:0]; // @[LZD.scala 49:47]
  assign _T_408 = _T_401[1:0]; // @[LZD.scala 49:59]
  assign _T_409 = _T_402 ? _T_407 : _T_408; // @[LZD.scala 49:35]
  assign _T_411 = {_T_404,_T_406,_T_409}; // @[Cat.scala 29:58]
  assign _T_412 = sumXor[2:0]; // @[LZD.scala 44:32]
  assign _T_413 = _T_412[2:1]; // @[LZD.scala 43:32]
  assign _T_414 = _T_413 != 2'h0; // @[LZD.scala 39:14]
  assign _T_415 = _T_413[1]; // @[LZD.scala 39:21]
  assign _T_416 = _T_413[0]; // @[LZD.scala 39:30]
  assign _T_417 = ~ _T_416; // @[LZD.scala 39:27]
  assign _T_418 = _T_415 | _T_417; // @[LZD.scala 39:25]
  assign _T_419 = {_T_414,_T_418}; // @[Cat.scala 29:58]
  assign _T_420 = _T_412[0:0]; // @[LZD.scala 44:32]
  assign _T_422 = _T_419[1]; // @[Shift.scala 12:21]
  assign _T_424 = _T_419[0:0]; // @[LZD.scala 55:32]
  assign _T_425 = _T_422 ? _T_424 : _T_420; // @[LZD.scala 55:20]
  assign _T_427 = _T_411[3]; // @[Shift.scala 12:21]
  assign _T_429 = {1'h1,_T_422,_T_425}; // @[Cat.scala 29:58]
  assign _T_430 = _T_411[2:0]; // @[LZD.scala 55:32]
  assign _T_431 = _T_427 ? _T_430 : _T_429; // @[LZD.scala 55:20]
  assign sumLZD = {_T_427,_T_431}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 128:24]
  assign _T_432 = signSumSig[9:0]; // @[PositFMA.scala 129:38]
  assign _T_433 = shiftValue < 4'ha; // @[Shift.scala 16:24]
  assign _T_435 = shiftValue[3]; // @[Shift.scala 12:21]
  assign _T_436 = _T_432[1:0]; // @[Shift.scala 64:52]
  assign _T_438 = {_T_436,8'h0}; // @[Cat.scala 29:58]
  assign _T_439 = _T_435 ? _T_438 : _T_432; // @[Shift.scala 64:27]
  assign _T_440 = shiftValue[2:0]; // @[Shift.scala 66:70]
  assign _T_441 = _T_440[2]; // @[Shift.scala 12:21]
  assign _T_442 = _T_439[5:0]; // @[Shift.scala 64:52]
  assign _T_444 = {_T_442,4'h0}; // @[Cat.scala 29:58]
  assign _T_445 = _T_441 ? _T_444 : _T_439; // @[Shift.scala 64:27]
  assign _T_446 = _T_440[1:0]; // @[Shift.scala 66:70]
  assign _T_447 = _T_446[1]; // @[Shift.scala 12:21]
  assign _T_448 = _T_445[7:0]; // @[Shift.scala 64:52]
  assign _T_450 = {_T_448,2'h0}; // @[Cat.scala 29:58]
  assign _T_451 = _T_447 ? _T_450 : _T_445; // @[Shift.scala 64:27]
  assign _T_452 = _T_446[0:0]; // @[Shift.scala 66:70]
  assign _T_454 = _T_451[8:0]; // @[Shift.scala 64:52]
  assign _T_455 = {_T_454,1'h0}; // @[Cat.scala 29:58]
  assign _T_456 = _T_452 ? _T_455 : _T_451; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_433 ? _T_456 : 10'h0; // @[Shift.scala 16:10]
  assign _T_458 = $signed(greaterScale) + $signed(5'sh2); // @[PositFMA.scala 132:36]
  assign _T_459 = $signed(_T_458); // @[PositFMA.scala 132:36]
  assign _T_460 = {1'h1,_T_427,_T_431}; // @[Cat.scala 29:58]
  assign _T_461 = $signed(_T_460); // @[PositFMA.scala 132:61]
  assign _T_463 = $signed(_T_459) + $signed(_T_461); // @[PositFMA.scala 132:42]
  assign sumScale = $signed(_T_463); // @[PositFMA.scala 132:42]
  assign sumFrac = normalFracTmp[9:6]; // @[PositFMA.scala 133:41]
  assign grsTmp = normalFracTmp[5:0]; // @[PositFMA.scala 136:41]
  assign _T_464 = grsTmp[5:4]; // @[PositFMA.scala 139:40]
  assign _T_465 = grsTmp[3:0]; // @[PositFMA.scala 139:56]
  assign _T_466 = _T_465 != 4'h0; // @[PositFMA.scala 139:60]
  assign underflow = $signed(sumScale) < $signed(-5'sh6); // @[PositFMA.scala 146:32]
  assign overflow = $signed(sumScale) > $signed(5'sh5); // @[PositFMA.scala 147:32]
  assign _T_467 = signSumSig != 12'h0; // @[PositFMA.scala 156:32]
  assign decF_isZero = ~ _T_467; // @[PositFMA.scala 156:20]
  assign _T_469 = underflow ? $signed(-5'sh6) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_470 = overflow ? $signed(5'sh5) : $signed(_T_469); // @[Mux.scala 87:16]
  assign _GEN_18 = _T_470[3:0]; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  assign decF_scale = $signed(_GEN_18); // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  assign _T_472 = decF_scale[3:3]; // @[convert.scala 49:36]
  assign _T_474 = ~ decF_scale; // @[convert.scala 50:36]
  assign _T_475 = $signed(_T_474); // @[convert.scala 50:36]
  assign _T_476 = _T_472 ? $signed(_T_475) : $signed(decF_scale); // @[convert.scala 50:28]
  assign _T_477 = _T_472 ^ sumSign; // @[convert.scala 51:31]
  assign _T_478 = ~ _T_477; // @[convert.scala 53:34]
  assign _T_481 = {_T_478,_T_477,sumFrac,_T_464,_T_466}; // @[Cat.scala 29:58]
  assign _T_482 = $unsigned(_T_476); // @[Shift.scala 39:17]
  assign _T_483 = _T_482 < 4'h9; // @[Shift.scala 39:24]
  assign _T_485 = _T_481[8:8]; // @[Shift.scala 90:30]
  assign _T_486 = _T_481[7:0]; // @[Shift.scala 90:48]
  assign _T_487 = _T_486 != 8'h0; // @[Shift.scala 90:57]
  assign _T_488 = _T_485 | _T_487; // @[Shift.scala 90:39]
  assign _T_489 = _T_482[3]; // @[Shift.scala 12:21]
  assign _T_490 = _T_481[8]; // @[Shift.scala 12:21]
  assign _T_492 = _T_490 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_493 = {_T_492,_T_488}; // @[Cat.scala 29:58]
  assign _T_494 = _T_489 ? _T_493 : _T_481; // @[Shift.scala 91:22]
  assign _T_495 = _T_482[2:0]; // @[Shift.scala 92:77]
  assign _T_496 = _T_494[8:4]; // @[Shift.scala 90:30]
  assign _T_497 = _T_494[3:0]; // @[Shift.scala 90:48]
  assign _T_498 = _T_497 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_19 = {{4'd0}, _T_498}; // @[Shift.scala 90:39]
  assign _T_499 = _T_496 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_500 = _T_495[2]; // @[Shift.scala 12:21]
  assign _T_501 = _T_494[8]; // @[Shift.scala 12:21]
  assign _T_503 = _T_501 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_504 = {_T_503,_T_499}; // @[Cat.scala 29:58]
  assign _T_505 = _T_500 ? _T_504 : _T_494; // @[Shift.scala 91:22]
  assign _T_506 = _T_495[1:0]; // @[Shift.scala 92:77]
  assign _T_507 = _T_505[8:2]; // @[Shift.scala 90:30]
  assign _T_508 = _T_505[1:0]; // @[Shift.scala 90:48]
  assign _T_509 = _T_508 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{6'd0}, _T_509}; // @[Shift.scala 90:39]
  assign _T_510 = _T_507 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_511 = _T_506[1]; // @[Shift.scala 12:21]
  assign _T_512 = _T_505[8]; // @[Shift.scala 12:21]
  assign _T_514 = _T_512 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_515 = {_T_514,_T_510}; // @[Cat.scala 29:58]
  assign _T_516 = _T_511 ? _T_515 : _T_505; // @[Shift.scala 91:22]
  assign _T_517 = _T_506[0:0]; // @[Shift.scala 92:77]
  assign _T_518 = _T_516[8:1]; // @[Shift.scala 90:30]
  assign _T_519 = _T_516[0:0]; // @[Shift.scala 90:48]
  assign _GEN_21 = {{7'd0}, _T_519}; // @[Shift.scala 90:39]
  assign _T_521 = _T_518 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_523 = _T_516[8]; // @[Shift.scala 12:21]
  assign _T_524 = {_T_523,_T_521}; // @[Cat.scala 29:58]
  assign _T_525 = _T_517 ? _T_524 : _T_516; // @[Shift.scala 91:22]
  assign _T_528 = _T_490 ? 9'h1ff : 9'h0; // @[Bitwise.scala 71:12]
  assign _T_529 = _T_483 ? _T_525 : _T_528; // @[Shift.scala 39:10]
  assign _T_530 = _T_529[3]; // @[convert.scala 55:31]
  assign _T_531 = _T_529[2]; // @[convert.scala 56:31]
  assign _T_532 = _T_529[1]; // @[convert.scala 57:31]
  assign _T_533 = _T_529[0]; // @[convert.scala 58:31]
  assign _T_534 = _T_529[8:3]; // @[convert.scala 59:69]
  assign _T_535 = _T_534 != 6'h0; // @[convert.scala 59:81]
  assign _T_536 = ~ _T_535; // @[convert.scala 59:50]
  assign _T_538 = _T_534 == 6'h3f; // @[convert.scala 60:81]
  assign _T_539 = _T_530 | _T_532; // @[convert.scala 61:44]
  assign _T_540 = _T_539 | _T_533; // @[convert.scala 61:52]
  assign _T_541 = _T_531 & _T_540; // @[convert.scala 61:36]
  assign _T_542 = ~ _T_538; // @[convert.scala 62:63]
  assign _T_543 = _T_542 & _T_541; // @[convert.scala 62:103]
  assign _T_544 = _T_536 | _T_543; // @[convert.scala 62:60]
  assign _GEN_22 = {{5'd0}, _T_544}; // @[convert.scala 63:56]
  assign _T_547 = _T_534 + _GEN_22; // @[convert.scala 63:56]
  assign _T_548 = {sumSign,_T_547}; // @[Cat.scala 29:58]
  assign io_F = _T_556; // @[PositFMA.scala 176:15]
  assign io_outValid = _T_552; // @[PositFMA.scala 175:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulSig_phase2 = _RAND_1[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_552 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_556 = _RAND_9[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      if (_T_204) begin
        if (_T_211) begin
          addFrac_phase2 <= _T_214;
        end else begin
          if (_T_206) begin
            addFrac_phase2 <= _T_209;
          end else begin
            addFrac_phase2 <= _T_203;
          end
        end
      end else begin
        addFrac_phase2 <= 4'h0;
      end
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_163;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_552 <= 1'h0;
    end else begin
      _T_552 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_556 <= 7'h40;
      end else begin
        if (decF_isZero) begin
          _T_556 <= 7'h0;
        end else begin
          _T_556 <= _T_548;
        end
      end
    end
  end
endmodule
