module Shifter9_5(
  input        clock,
  input        reset,
  input  [8:0] io_in,
  input  [4:0] io_shiftamt,
  output [8:0] io_shiftout
);
  wire  _T; // @[Shift.scala 39:24]
  wire [3:0] _T_1; // @[Shift.scala 40:44]
  wire  _T_2; // @[Shift.scala 90:30]
  wire [7:0] _T_3; // @[Shift.scala 90:48]
  wire  _T_4; // @[Shift.scala 90:57]
  wire  _T_5; // @[Shift.scala 90:39]
  wire  _T_6; // @[Shift.scala 12:21]
  wire  _T_7; // @[Shift.scala 12:21]
  wire [7:0] _T_9; // @[Bitwise.scala 71:12]
  wire [8:0] _T_10; // @[Cat.scala 29:58]
  wire [8:0] _T_11; // @[Shift.scala 91:22]
  wire [2:0] _T_12; // @[Shift.scala 92:77]
  wire [4:0] _T_13; // @[Shift.scala 90:30]
  wire [3:0] _T_14; // @[Shift.scala 90:48]
  wire  _T_15; // @[Shift.scala 90:57]
  wire [4:0] _GEN_0; // @[Shift.scala 90:39]
  wire [4:0] _T_16; // @[Shift.scala 90:39]
  wire  _T_17; // @[Shift.scala 12:21]
  wire  _T_18; // @[Shift.scala 12:21]
  wire [3:0] _T_20; // @[Bitwise.scala 71:12]
  wire [8:0] _T_21; // @[Cat.scala 29:58]
  wire [8:0] _T_22; // @[Shift.scala 91:22]
  wire [1:0] _T_23; // @[Shift.scala 92:77]
  wire [6:0] _T_24; // @[Shift.scala 90:30]
  wire [1:0] _T_25; // @[Shift.scala 90:48]
  wire  _T_26; // @[Shift.scala 90:57]
  wire [6:0] _GEN_1; // @[Shift.scala 90:39]
  wire [6:0] _T_27; // @[Shift.scala 90:39]
  wire  _T_28; // @[Shift.scala 12:21]
  wire  _T_29; // @[Shift.scala 12:21]
  wire [1:0] _T_31; // @[Bitwise.scala 71:12]
  wire [8:0] _T_32; // @[Cat.scala 29:58]
  wire [8:0] _T_33; // @[Shift.scala 91:22]
  wire  _T_34; // @[Shift.scala 92:77]
  wire [7:0] _T_35; // @[Shift.scala 90:30]
  wire  _T_36; // @[Shift.scala 90:48]
  wire [7:0] _GEN_2; // @[Shift.scala 90:39]
  wire [7:0] _T_38; // @[Shift.scala 90:39]
  wire  _T_40; // @[Shift.scala 12:21]
  wire [8:0] _T_41; // @[Cat.scala 29:58]
  wire [8:0] _T_42; // @[Shift.scala 91:22]
  wire [8:0] _T_45; // @[Bitwise.scala 71:12]
  assign _T = io_shiftamt < 5'h9; // @[Shift.scala 39:24]
  assign _T_1 = io_shiftamt[3:0]; // @[Shift.scala 40:44]
  assign _T_2 = io_in[8:8]; // @[Shift.scala 90:30]
  assign _T_3 = io_in[7:0]; // @[Shift.scala 90:48]
  assign _T_4 = _T_3 != 8'h0; // @[Shift.scala 90:57]
  assign _T_5 = _T_2 | _T_4; // @[Shift.scala 90:39]
  assign _T_6 = _T_1[3]; // @[Shift.scala 12:21]
  assign _T_7 = io_in[8]; // @[Shift.scala 12:21]
  assign _T_9 = _T_7 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_10 = {_T_9,_T_5}; // @[Cat.scala 29:58]
  assign _T_11 = _T_6 ? _T_10 : io_in; // @[Shift.scala 91:22]
  assign _T_12 = _T_1[2:0]; // @[Shift.scala 92:77]
  assign _T_13 = _T_11[8:4]; // @[Shift.scala 90:30]
  assign _T_14 = _T_11[3:0]; // @[Shift.scala 90:48]
  assign _T_15 = _T_14 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{4'd0}, _T_15}; // @[Shift.scala 90:39]
  assign _T_16 = _T_13 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_17 = _T_12[2]; // @[Shift.scala 12:21]
  assign _T_18 = _T_11[8]; // @[Shift.scala 12:21]
  assign _T_20 = _T_18 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_21 = {_T_20,_T_16}; // @[Cat.scala 29:58]
  assign _T_22 = _T_17 ? _T_21 : _T_11; // @[Shift.scala 91:22]
  assign _T_23 = _T_12[1:0]; // @[Shift.scala 92:77]
  assign _T_24 = _T_22[8:2]; // @[Shift.scala 90:30]
  assign _T_25 = _T_22[1:0]; // @[Shift.scala 90:48]
  assign _T_26 = _T_25 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{6'd0}, _T_26}; // @[Shift.scala 90:39]
  assign _T_27 = _T_24 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_28 = _T_23[1]; // @[Shift.scala 12:21]
  assign _T_29 = _T_22[8]; // @[Shift.scala 12:21]
  assign _T_31 = _T_29 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_32 = {_T_31,_T_27}; // @[Cat.scala 29:58]
  assign _T_33 = _T_28 ? _T_32 : _T_22; // @[Shift.scala 91:22]
  assign _T_34 = _T_23[0:0]; // @[Shift.scala 92:77]
  assign _T_35 = _T_33[8:1]; // @[Shift.scala 90:30]
  assign _T_36 = _T_33[0:0]; // @[Shift.scala 90:48]
  assign _GEN_2 = {{7'd0}, _T_36}; // @[Shift.scala 90:39]
  assign _T_38 = _T_35 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_40 = _T_33[8]; // @[Shift.scala 12:21]
  assign _T_41 = {_T_40,_T_38}; // @[Cat.scala 29:58]
  assign _T_42 = _T_34 ? _T_41 : _T_33; // @[Shift.scala 91:22]
  assign _T_45 = _T_7 ? 9'h1ff : 9'h0; // @[Bitwise.scala 71:12]
  assign io_shiftout = _T ? _T_42 : _T_45; // @[Shif.scala 16:15]
endmodule
