module QuireToPosit6_8_0(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [31:0] io_quireIn,
  output [7:0]  io_positOut,
  output        io_outValid
);
  wire [30:0] _T; // @[QuireToPosit.scala 47:43]
  wire  _T_1; // @[QuireToPosit.scala 47:47]
  wire  tailIsZero; // @[QuireToPosit.scala 47:27]
  wire  _T_2; // @[QuireToPosit.scala 49:45]
  wire  outRawFloat_isNaR; // @[QuireToPosit.scala 49:49]
  wire  _T_5; // @[QuireToPosit.scala 50:31]
  wire  outRawFloat_isZero; // @[QuireToPosit.scala 50:51]
  wire [30:0] _T_8; // @[QuireToPosit.scala 58:41]
  wire [30:0] _T_9; // @[QuireToPosit.scala 58:68]
  wire [30:0] quireXOR; // @[QuireToPosit.scala 58:56]
  wire [15:0] _T_10; // @[LZD.scala 43:32]
  wire [7:0] _T_11; // @[LZD.scala 43:32]
  wire [3:0] _T_12; // @[LZD.scala 43:32]
  wire [1:0] _T_13; // @[LZD.scala 43:32]
  wire  _T_14; // @[LZD.scala 39:14]
  wire  _T_15; // @[LZD.scala 39:21]
  wire  _T_16; // @[LZD.scala 39:30]
  wire  _T_17; // @[LZD.scala 39:27]
  wire  _T_18; // @[LZD.scala 39:25]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire [1:0] _T_20; // @[LZD.scala 44:32]
  wire  _T_21; // @[LZD.scala 39:14]
  wire  _T_22; // @[LZD.scala 39:21]
  wire  _T_23; // @[LZD.scala 39:30]
  wire  _T_24; // @[LZD.scala 39:27]
  wire  _T_25; // @[LZD.scala 39:25]
  wire [1:0] _T_26; // @[Cat.scala 29:58]
  wire  _T_27; // @[Shift.scala 12:21]
  wire  _T_28; // @[Shift.scala 12:21]
  wire  _T_29; // @[LZD.scala 49:16]
  wire  _T_30; // @[LZD.scala 49:27]
  wire  _T_31; // @[LZD.scala 49:25]
  wire  _T_32; // @[LZD.scala 49:47]
  wire  _T_33; // @[LZD.scala 49:59]
  wire  _T_34; // @[LZD.scala 49:35]
  wire [2:0] _T_36; // @[Cat.scala 29:58]
  wire [3:0] _T_37; // @[LZD.scala 44:32]
  wire [1:0] _T_38; // @[LZD.scala 43:32]
  wire  _T_39; // @[LZD.scala 39:14]
  wire  _T_40; // @[LZD.scala 39:21]
  wire  _T_41; // @[LZD.scala 39:30]
  wire  _T_42; // @[LZD.scala 39:27]
  wire  _T_43; // @[LZD.scala 39:25]
  wire [1:0] _T_44; // @[Cat.scala 29:58]
  wire [1:0] _T_45; // @[LZD.scala 44:32]
  wire  _T_46; // @[LZD.scala 39:14]
  wire  _T_47; // @[LZD.scala 39:21]
  wire  _T_48; // @[LZD.scala 39:30]
  wire  _T_49; // @[LZD.scala 39:27]
  wire  _T_50; // @[LZD.scala 39:25]
  wire [1:0] _T_51; // @[Cat.scala 29:58]
  wire  _T_52; // @[Shift.scala 12:21]
  wire  _T_53; // @[Shift.scala 12:21]
  wire  _T_54; // @[LZD.scala 49:16]
  wire  _T_55; // @[LZD.scala 49:27]
  wire  _T_56; // @[LZD.scala 49:25]
  wire  _T_57; // @[LZD.scala 49:47]
  wire  _T_58; // @[LZD.scala 49:59]
  wire  _T_59; // @[LZD.scala 49:35]
  wire [2:0] _T_61; // @[Cat.scala 29:58]
  wire  _T_62; // @[Shift.scala 12:21]
  wire  _T_63; // @[Shift.scala 12:21]
  wire  _T_64; // @[LZD.scala 49:16]
  wire  _T_65; // @[LZD.scala 49:27]
  wire  _T_66; // @[LZD.scala 49:25]
  wire [1:0] _T_67; // @[LZD.scala 49:47]
  wire [1:0] _T_68; // @[LZD.scala 49:59]
  wire [1:0] _T_69; // @[LZD.scala 49:35]
  wire [3:0] _T_71; // @[Cat.scala 29:58]
  wire [7:0] _T_72; // @[LZD.scala 44:32]
  wire [3:0] _T_73; // @[LZD.scala 43:32]
  wire [1:0] _T_74; // @[LZD.scala 43:32]
  wire  _T_75; // @[LZD.scala 39:14]
  wire  _T_76; // @[LZD.scala 39:21]
  wire  _T_77; // @[LZD.scala 39:30]
  wire  _T_78; // @[LZD.scala 39:27]
  wire  _T_79; // @[LZD.scala 39:25]
  wire [1:0] _T_80; // @[Cat.scala 29:58]
  wire [1:0] _T_81; // @[LZD.scala 44:32]
  wire  _T_82; // @[LZD.scala 39:14]
  wire  _T_83; // @[LZD.scala 39:21]
  wire  _T_84; // @[LZD.scala 39:30]
  wire  _T_85; // @[LZD.scala 39:27]
  wire  _T_86; // @[LZD.scala 39:25]
  wire [1:0] _T_87; // @[Cat.scala 29:58]
  wire  _T_88; // @[Shift.scala 12:21]
  wire  _T_89; // @[Shift.scala 12:21]
  wire  _T_90; // @[LZD.scala 49:16]
  wire  _T_91; // @[LZD.scala 49:27]
  wire  _T_92; // @[LZD.scala 49:25]
  wire  _T_93; // @[LZD.scala 49:47]
  wire  _T_94; // @[LZD.scala 49:59]
  wire  _T_95; // @[LZD.scala 49:35]
  wire [2:0] _T_97; // @[Cat.scala 29:58]
  wire [3:0] _T_98; // @[LZD.scala 44:32]
  wire [1:0] _T_99; // @[LZD.scala 43:32]
  wire  _T_100; // @[LZD.scala 39:14]
  wire  _T_101; // @[LZD.scala 39:21]
  wire  _T_102; // @[LZD.scala 39:30]
  wire  _T_103; // @[LZD.scala 39:27]
  wire  _T_104; // @[LZD.scala 39:25]
  wire [1:0] _T_105; // @[Cat.scala 29:58]
  wire [1:0] _T_106; // @[LZD.scala 44:32]
  wire  _T_107; // @[LZD.scala 39:14]
  wire  _T_108; // @[LZD.scala 39:21]
  wire  _T_109; // @[LZD.scala 39:30]
  wire  _T_110; // @[LZD.scala 39:27]
  wire  _T_111; // @[LZD.scala 39:25]
  wire [1:0] _T_112; // @[Cat.scala 29:58]
  wire  _T_113; // @[Shift.scala 12:21]
  wire  _T_114; // @[Shift.scala 12:21]
  wire  _T_115; // @[LZD.scala 49:16]
  wire  _T_116; // @[LZD.scala 49:27]
  wire  _T_117; // @[LZD.scala 49:25]
  wire  _T_118; // @[LZD.scala 49:47]
  wire  _T_119; // @[LZD.scala 49:59]
  wire  _T_120; // @[LZD.scala 49:35]
  wire [2:0] _T_122; // @[Cat.scala 29:58]
  wire  _T_123; // @[Shift.scala 12:21]
  wire  _T_124; // @[Shift.scala 12:21]
  wire  _T_125; // @[LZD.scala 49:16]
  wire  _T_126; // @[LZD.scala 49:27]
  wire  _T_127; // @[LZD.scala 49:25]
  wire [1:0] _T_128; // @[LZD.scala 49:47]
  wire [1:0] _T_129; // @[LZD.scala 49:59]
  wire [1:0] _T_130; // @[LZD.scala 49:35]
  wire [3:0] _T_132; // @[Cat.scala 29:58]
  wire  _T_133; // @[Shift.scala 12:21]
  wire  _T_134; // @[Shift.scala 12:21]
  wire  _T_135; // @[LZD.scala 49:16]
  wire  _T_136; // @[LZD.scala 49:27]
  wire  _T_137; // @[LZD.scala 49:25]
  wire [2:0] _T_138; // @[LZD.scala 49:47]
  wire [2:0] _T_139; // @[LZD.scala 49:59]
  wire [2:0] _T_140; // @[LZD.scala 49:35]
  wire [4:0] _T_142; // @[Cat.scala 29:58]
  wire [14:0] _T_143; // @[LZD.scala 44:32]
  wire [7:0] _T_144; // @[LZD.scala 43:32]
  wire [3:0] _T_145; // @[LZD.scala 43:32]
  wire [1:0] _T_146; // @[LZD.scala 43:32]
  wire  _T_147; // @[LZD.scala 39:14]
  wire  _T_148; // @[LZD.scala 39:21]
  wire  _T_149; // @[LZD.scala 39:30]
  wire  _T_150; // @[LZD.scala 39:27]
  wire  _T_151; // @[LZD.scala 39:25]
  wire [1:0] _T_152; // @[Cat.scala 29:58]
  wire [1:0] _T_153; // @[LZD.scala 44:32]
  wire  _T_154; // @[LZD.scala 39:14]
  wire  _T_155; // @[LZD.scala 39:21]
  wire  _T_156; // @[LZD.scala 39:30]
  wire  _T_157; // @[LZD.scala 39:27]
  wire  _T_158; // @[LZD.scala 39:25]
  wire [1:0] _T_159; // @[Cat.scala 29:58]
  wire  _T_160; // @[Shift.scala 12:21]
  wire  _T_161; // @[Shift.scala 12:21]
  wire  _T_162; // @[LZD.scala 49:16]
  wire  _T_163; // @[LZD.scala 49:27]
  wire  _T_164; // @[LZD.scala 49:25]
  wire  _T_165; // @[LZD.scala 49:47]
  wire  _T_166; // @[LZD.scala 49:59]
  wire  _T_167; // @[LZD.scala 49:35]
  wire [2:0] _T_169; // @[Cat.scala 29:58]
  wire [3:0] _T_170; // @[LZD.scala 44:32]
  wire [1:0] _T_171; // @[LZD.scala 43:32]
  wire  _T_172; // @[LZD.scala 39:14]
  wire  _T_173; // @[LZD.scala 39:21]
  wire  _T_174; // @[LZD.scala 39:30]
  wire  _T_175; // @[LZD.scala 39:27]
  wire  _T_176; // @[LZD.scala 39:25]
  wire [1:0] _T_177; // @[Cat.scala 29:58]
  wire [1:0] _T_178; // @[LZD.scala 44:32]
  wire  _T_179; // @[LZD.scala 39:14]
  wire  _T_180; // @[LZD.scala 39:21]
  wire  _T_181; // @[LZD.scala 39:30]
  wire  _T_182; // @[LZD.scala 39:27]
  wire  _T_183; // @[LZD.scala 39:25]
  wire [1:0] _T_184; // @[Cat.scala 29:58]
  wire  _T_185; // @[Shift.scala 12:21]
  wire  _T_186; // @[Shift.scala 12:21]
  wire  _T_187; // @[LZD.scala 49:16]
  wire  _T_188; // @[LZD.scala 49:27]
  wire  _T_189; // @[LZD.scala 49:25]
  wire  _T_190; // @[LZD.scala 49:47]
  wire  _T_191; // @[LZD.scala 49:59]
  wire  _T_192; // @[LZD.scala 49:35]
  wire [2:0] _T_194; // @[Cat.scala 29:58]
  wire  _T_195; // @[Shift.scala 12:21]
  wire  _T_196; // @[Shift.scala 12:21]
  wire  _T_197; // @[LZD.scala 49:16]
  wire  _T_198; // @[LZD.scala 49:27]
  wire  _T_199; // @[LZD.scala 49:25]
  wire [1:0] _T_200; // @[LZD.scala 49:47]
  wire [1:0] _T_201; // @[LZD.scala 49:59]
  wire [1:0] _T_202; // @[LZD.scala 49:35]
  wire [3:0] _T_204; // @[Cat.scala 29:58]
  wire [6:0] _T_205; // @[LZD.scala 44:32]
  wire [3:0] _T_206; // @[LZD.scala 43:32]
  wire [1:0] _T_207; // @[LZD.scala 43:32]
  wire  _T_208; // @[LZD.scala 39:14]
  wire  _T_209; // @[LZD.scala 39:21]
  wire  _T_210; // @[LZD.scala 39:30]
  wire  _T_211; // @[LZD.scala 39:27]
  wire  _T_212; // @[LZD.scala 39:25]
  wire [1:0] _T_213; // @[Cat.scala 29:58]
  wire [1:0] _T_214; // @[LZD.scala 44:32]
  wire  _T_215; // @[LZD.scala 39:14]
  wire  _T_216; // @[LZD.scala 39:21]
  wire  _T_217; // @[LZD.scala 39:30]
  wire  _T_218; // @[LZD.scala 39:27]
  wire  _T_219; // @[LZD.scala 39:25]
  wire [1:0] _T_220; // @[Cat.scala 29:58]
  wire  _T_221; // @[Shift.scala 12:21]
  wire  _T_222; // @[Shift.scala 12:21]
  wire  _T_223; // @[LZD.scala 49:16]
  wire  _T_224; // @[LZD.scala 49:27]
  wire  _T_225; // @[LZD.scala 49:25]
  wire  _T_226; // @[LZD.scala 49:47]
  wire  _T_227; // @[LZD.scala 49:59]
  wire  _T_228; // @[LZD.scala 49:35]
  wire [2:0] _T_230; // @[Cat.scala 29:58]
  wire [2:0] _T_231; // @[LZD.scala 44:32]
  wire [1:0] _T_232; // @[LZD.scala 43:32]
  wire  _T_233; // @[LZD.scala 39:14]
  wire  _T_234; // @[LZD.scala 39:21]
  wire  _T_235; // @[LZD.scala 39:30]
  wire  _T_236; // @[LZD.scala 39:27]
  wire  _T_237; // @[LZD.scala 39:25]
  wire [1:0] _T_238; // @[Cat.scala 29:58]
  wire  _T_239; // @[LZD.scala 44:32]
  wire  _T_241; // @[Shift.scala 12:21]
  wire  _T_243; // @[LZD.scala 55:32]
  wire  _T_244; // @[LZD.scala 55:20]
  wire [1:0] _T_245; // @[Cat.scala 29:58]
  wire  _T_246; // @[Shift.scala 12:21]
  wire [1:0] _T_248; // @[LZD.scala 55:32]
  wire [1:0] _T_249; // @[LZD.scala 55:20]
  wire [2:0] _T_250; // @[Cat.scala 29:58]
  wire  _T_251; // @[Shift.scala 12:21]
  wire [2:0] _T_253; // @[LZD.scala 55:32]
  wire [2:0] _T_254; // @[LZD.scala 55:20]
  wire [3:0] _T_255; // @[Cat.scala 29:58]
  wire  _T_256; // @[Shift.scala 12:21]
  wire [3:0] _T_258; // @[LZD.scala 55:32]
  wire [3:0] _T_259; // @[LZD.scala 55:20]
  wire [5:0] scaleBias; // @[Cat.scala 29:58]
  wire [5:0] _T_260; // @[QuireToPosit.scala 61:53]
  wire [6:0] _GEN_2; // @[QuireToPosit.scala 61:41]
  wire [6:0] _T_262; // @[QuireToPosit.scala 61:41]
  wire [6:0] realScale; // @[QuireToPosit.scala 61:41]
  wire  underflow; // @[QuireToPosit.scala 62:41]
  wire  overflow; // @[QuireToPosit.scala 63:35]
  wire [6:0] _T_263; // @[Mux.scala 87:16]
  wire [6:0] _T_264; // @[Mux.scala 87:16]
  wire  _T_265; // @[Abs.scala 10:21]
  wire [6:0] _T_267; // @[Bitwise.scala 71:12]
  wire [6:0] _T_268; // @[Abs.scala 10:31]
  wire [6:0] _T_269; // @[Abs.scala 10:26]
  wire [6:0] _GEN_3; // @[Abs.scala 10:39]
  wire [6:0] absRealScale; // @[Abs.scala 10:39]
  wire  _T_272; // @[Shift.scala 16:24]
  wire [4:0] _T_273; // @[Shift.scala 17:37]
  wire  _T_274; // @[Shift.scala 12:21]
  wire [15:0] _T_275; // @[Shift.scala 64:52]
  wire [31:0] _T_277; // @[Cat.scala 29:58]
  wire [31:0] _T_278; // @[Shift.scala 64:27]
  wire [3:0] _T_279; // @[Shift.scala 66:70]
  wire  _T_280; // @[Shift.scala 12:21]
  wire [23:0] _T_281; // @[Shift.scala 64:52]
  wire [31:0] _T_283; // @[Cat.scala 29:58]
  wire [31:0] _T_284; // @[Shift.scala 64:27]
  wire [2:0] _T_285; // @[Shift.scala 66:70]
  wire  _T_286; // @[Shift.scala 12:21]
  wire [27:0] _T_287; // @[Shift.scala 64:52]
  wire [31:0] _T_289; // @[Cat.scala 29:58]
  wire [31:0] _T_290; // @[Shift.scala 64:27]
  wire [1:0] _T_291; // @[Shift.scala 66:70]
  wire  _T_292; // @[Shift.scala 12:21]
  wire [29:0] _T_293; // @[Shift.scala 64:52]
  wire [31:0] _T_295; // @[Cat.scala 29:58]
  wire [31:0] _T_296; // @[Shift.scala 64:27]
  wire  _T_297; // @[Shift.scala 66:70]
  wire [30:0] _T_299; // @[Shift.scala 64:52]
  wire [31:0] _T_300; // @[Cat.scala 29:58]
  wire [31:0] _T_301; // @[Shift.scala 64:27]
  wire [31:0] quireLeftShift; // @[Shift.scala 16:10]
  wire [15:0] _T_306; // @[Shift.scala 77:66]
  wire [31:0] _T_307; // @[Cat.scala 29:58]
  wire [31:0] _T_308; // @[Shift.scala 77:22]
  wire [23:0] _T_312; // @[Shift.scala 77:66]
  wire [31:0] _T_313; // @[Cat.scala 29:58]
  wire [31:0] _T_314; // @[Shift.scala 77:22]
  wire [27:0] _T_318; // @[Shift.scala 77:66]
  wire [31:0] _T_319; // @[Cat.scala 29:58]
  wire [31:0] _T_320; // @[Shift.scala 77:22]
  wire [29:0] _T_324; // @[Shift.scala 77:66]
  wire [31:0] _T_325; // @[Cat.scala 29:58]
  wire [31:0] _T_326; // @[Shift.scala 77:22]
  wire [30:0] _T_329; // @[Shift.scala 77:66]
  wire [31:0] _T_330; // @[Cat.scala 29:58]
  wire [31:0] _T_331; // @[Shift.scala 77:22]
  wire [31:0] quireRightShift; // @[Shift.scala 27:10]
  wire [6:0] _T_333; // @[QuireToPosit.scala 89:49]
  wire [4:0] _T_334; // @[QuireToPosit.scala 90:127]
  wire  _T_335; // @[QuireToPosit.scala 90:154]
  wire [7:0] realFGRSTmp1; // @[Cat.scala 29:58]
  wire [6:0] _T_336; // @[QuireToPosit.scala 91:50]
  wire [4:0] _T_337; // @[QuireToPosit.scala 92:128]
  wire  _T_338; // @[QuireToPosit.scala 92:155]
  wire [7:0] realFGRSTmp2; // @[Cat.scala 29:58]
  wire [7:0] realFGRS; // @[QuireToPosit.scala 93:34]
  wire [4:0] outRawFloat_fraction; // @[QuireToPosit.scala 95:46]
  wire [2:0] outRawFloat_grs; // @[QuireToPosit.scala 96:46]
  wire [3:0] _GEN_4; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  wire [3:0] outRawFloat_scale; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  wire  _T_344; // @[convert.scala 49:36]
  wire [3:0] _T_346; // @[convert.scala 50:36]
  wire [3:0] _T_347; // @[convert.scala 50:36]
  wire [3:0] _T_348; // @[convert.scala 50:28]
  wire  _T_349; // @[convert.scala 51:31]
  wire  _T_350; // @[convert.scala 53:34]
  wire [9:0] _T_353; // @[Cat.scala 29:58]
  wire [3:0] _T_354; // @[Shift.scala 39:17]
  wire  _T_355; // @[Shift.scala 39:24]
  wire [1:0] _T_357; // @[Shift.scala 90:30]
  wire [7:0] _T_358; // @[Shift.scala 90:48]
  wire  _T_359; // @[Shift.scala 90:57]
  wire [1:0] _GEN_5; // @[Shift.scala 90:39]
  wire [1:0] _T_360; // @[Shift.scala 90:39]
  wire  _T_361; // @[Shift.scala 12:21]
  wire  _T_362; // @[Shift.scala 12:21]
  wire [7:0] _T_364; // @[Bitwise.scala 71:12]
  wire [9:0] _T_365; // @[Cat.scala 29:58]
  wire [9:0] _T_366; // @[Shift.scala 91:22]
  wire [2:0] _T_367; // @[Shift.scala 92:77]
  wire [5:0] _T_368; // @[Shift.scala 90:30]
  wire [3:0] _T_369; // @[Shift.scala 90:48]
  wire  _T_370; // @[Shift.scala 90:57]
  wire [5:0] _GEN_6; // @[Shift.scala 90:39]
  wire [5:0] _T_371; // @[Shift.scala 90:39]
  wire  _T_372; // @[Shift.scala 12:21]
  wire  _T_373; // @[Shift.scala 12:21]
  wire [3:0] _T_375; // @[Bitwise.scala 71:12]
  wire [9:0] _T_376; // @[Cat.scala 29:58]
  wire [9:0] _T_377; // @[Shift.scala 91:22]
  wire [1:0] _T_378; // @[Shift.scala 92:77]
  wire [7:0] _T_379; // @[Shift.scala 90:30]
  wire [1:0] _T_380; // @[Shift.scala 90:48]
  wire  _T_381; // @[Shift.scala 90:57]
  wire [7:0] _GEN_7; // @[Shift.scala 90:39]
  wire [7:0] _T_382; // @[Shift.scala 90:39]
  wire  _T_383; // @[Shift.scala 12:21]
  wire  _T_384; // @[Shift.scala 12:21]
  wire [1:0] _T_386; // @[Bitwise.scala 71:12]
  wire [9:0] _T_387; // @[Cat.scala 29:58]
  wire [9:0] _T_388; // @[Shift.scala 91:22]
  wire  _T_389; // @[Shift.scala 92:77]
  wire [8:0] _T_390; // @[Shift.scala 90:30]
  wire  _T_391; // @[Shift.scala 90:48]
  wire [8:0] _GEN_8; // @[Shift.scala 90:39]
  wire [8:0] _T_393; // @[Shift.scala 90:39]
  wire  _T_395; // @[Shift.scala 12:21]
  wire [9:0] _T_396; // @[Cat.scala 29:58]
  wire [9:0] _T_397; // @[Shift.scala 91:22]
  wire [9:0] _T_400; // @[Bitwise.scala 71:12]
  wire [9:0] _T_401; // @[Shift.scala 39:10]
  wire  _T_402; // @[convert.scala 55:31]
  wire  _T_403; // @[convert.scala 56:31]
  wire  _T_404; // @[convert.scala 57:31]
  wire  _T_405; // @[convert.scala 58:31]
  wire [6:0] _T_406; // @[convert.scala 59:69]
  wire  _T_407; // @[convert.scala 59:81]
  wire  _T_408; // @[convert.scala 59:50]
  wire  _T_410; // @[convert.scala 60:81]
  wire  _T_411; // @[convert.scala 61:44]
  wire  _T_412; // @[convert.scala 61:52]
  wire  _T_413; // @[convert.scala 61:36]
  wire  _T_414; // @[convert.scala 62:63]
  wire  _T_415; // @[convert.scala 62:103]
  wire  _T_416; // @[convert.scala 62:60]
  wire [6:0] _GEN_9; // @[convert.scala 63:56]
  wire [6:0] _T_419; // @[convert.scala 63:56]
  wire [7:0] _T_420; // @[Cat.scala 29:58]
  reg  _T_424; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [7:0] _T_428; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  assign _T = io_quireIn[30:0]; // @[QuireToPosit.scala 47:43]
  assign _T_1 = _T != 31'h0; // @[QuireToPosit.scala 47:47]
  assign tailIsZero = ~ _T_1; // @[QuireToPosit.scala 47:27]
  assign _T_2 = io_quireIn[31:31]; // @[QuireToPosit.scala 49:45]
  assign outRawFloat_isNaR = _T_2 & tailIsZero; // @[QuireToPosit.scala 49:49]
  assign _T_5 = ~ _T_2; // @[QuireToPosit.scala 50:31]
  assign outRawFloat_isZero = _T_5 & tailIsZero; // @[QuireToPosit.scala 50:51]
  assign _T_8 = io_quireIn[31:1]; // @[QuireToPosit.scala 58:41]
  assign _T_9 = io_quireIn[30:0]; // @[QuireToPosit.scala 58:68]
  assign quireXOR = _T_8 ^ _T_9; // @[QuireToPosit.scala 58:56]
  assign _T_10 = quireXOR[30:15]; // @[LZD.scala 43:32]
  assign _T_11 = _T_10[15:8]; // @[LZD.scala 43:32]
  assign _T_12 = _T_11[7:4]; // @[LZD.scala 43:32]
  assign _T_13 = _T_12[3:2]; // @[LZD.scala 43:32]
  assign _T_14 = _T_13 != 2'h0; // @[LZD.scala 39:14]
  assign _T_15 = _T_13[1]; // @[LZD.scala 39:21]
  assign _T_16 = _T_13[0]; // @[LZD.scala 39:30]
  assign _T_17 = ~ _T_16; // @[LZD.scala 39:27]
  assign _T_18 = _T_15 | _T_17; // @[LZD.scala 39:25]
  assign _T_19 = {_T_14,_T_18}; // @[Cat.scala 29:58]
  assign _T_20 = _T_12[1:0]; // @[LZD.scala 44:32]
  assign _T_21 = _T_20 != 2'h0; // @[LZD.scala 39:14]
  assign _T_22 = _T_20[1]; // @[LZD.scala 39:21]
  assign _T_23 = _T_20[0]; // @[LZD.scala 39:30]
  assign _T_24 = ~ _T_23; // @[LZD.scala 39:27]
  assign _T_25 = _T_22 | _T_24; // @[LZD.scala 39:25]
  assign _T_26 = {_T_21,_T_25}; // @[Cat.scala 29:58]
  assign _T_27 = _T_19[1]; // @[Shift.scala 12:21]
  assign _T_28 = _T_26[1]; // @[Shift.scala 12:21]
  assign _T_29 = _T_27 | _T_28; // @[LZD.scala 49:16]
  assign _T_30 = ~ _T_28; // @[LZD.scala 49:27]
  assign _T_31 = _T_27 | _T_30; // @[LZD.scala 49:25]
  assign _T_32 = _T_19[0:0]; // @[LZD.scala 49:47]
  assign _T_33 = _T_26[0:0]; // @[LZD.scala 49:59]
  assign _T_34 = _T_27 ? _T_32 : _T_33; // @[LZD.scala 49:35]
  assign _T_36 = {_T_29,_T_31,_T_34}; // @[Cat.scala 29:58]
  assign _T_37 = _T_11[3:0]; // @[LZD.scala 44:32]
  assign _T_38 = _T_37[3:2]; // @[LZD.scala 43:32]
  assign _T_39 = _T_38 != 2'h0; // @[LZD.scala 39:14]
  assign _T_40 = _T_38[1]; // @[LZD.scala 39:21]
  assign _T_41 = _T_38[0]; // @[LZD.scala 39:30]
  assign _T_42 = ~ _T_41; // @[LZD.scala 39:27]
  assign _T_43 = _T_40 | _T_42; // @[LZD.scala 39:25]
  assign _T_44 = {_T_39,_T_43}; // @[Cat.scala 29:58]
  assign _T_45 = _T_37[1:0]; // @[LZD.scala 44:32]
  assign _T_46 = _T_45 != 2'h0; // @[LZD.scala 39:14]
  assign _T_47 = _T_45[1]; // @[LZD.scala 39:21]
  assign _T_48 = _T_45[0]; // @[LZD.scala 39:30]
  assign _T_49 = ~ _T_48; // @[LZD.scala 39:27]
  assign _T_50 = _T_47 | _T_49; // @[LZD.scala 39:25]
  assign _T_51 = {_T_46,_T_50}; // @[Cat.scala 29:58]
  assign _T_52 = _T_44[1]; // @[Shift.scala 12:21]
  assign _T_53 = _T_51[1]; // @[Shift.scala 12:21]
  assign _T_54 = _T_52 | _T_53; // @[LZD.scala 49:16]
  assign _T_55 = ~ _T_53; // @[LZD.scala 49:27]
  assign _T_56 = _T_52 | _T_55; // @[LZD.scala 49:25]
  assign _T_57 = _T_44[0:0]; // @[LZD.scala 49:47]
  assign _T_58 = _T_51[0:0]; // @[LZD.scala 49:59]
  assign _T_59 = _T_52 ? _T_57 : _T_58; // @[LZD.scala 49:35]
  assign _T_61 = {_T_54,_T_56,_T_59}; // @[Cat.scala 29:58]
  assign _T_62 = _T_36[2]; // @[Shift.scala 12:21]
  assign _T_63 = _T_61[2]; // @[Shift.scala 12:21]
  assign _T_64 = _T_62 | _T_63; // @[LZD.scala 49:16]
  assign _T_65 = ~ _T_63; // @[LZD.scala 49:27]
  assign _T_66 = _T_62 | _T_65; // @[LZD.scala 49:25]
  assign _T_67 = _T_36[1:0]; // @[LZD.scala 49:47]
  assign _T_68 = _T_61[1:0]; // @[LZD.scala 49:59]
  assign _T_69 = _T_62 ? _T_67 : _T_68; // @[LZD.scala 49:35]
  assign _T_71 = {_T_64,_T_66,_T_69}; // @[Cat.scala 29:58]
  assign _T_72 = _T_10[7:0]; // @[LZD.scala 44:32]
  assign _T_73 = _T_72[7:4]; // @[LZD.scala 43:32]
  assign _T_74 = _T_73[3:2]; // @[LZD.scala 43:32]
  assign _T_75 = _T_74 != 2'h0; // @[LZD.scala 39:14]
  assign _T_76 = _T_74[1]; // @[LZD.scala 39:21]
  assign _T_77 = _T_74[0]; // @[LZD.scala 39:30]
  assign _T_78 = ~ _T_77; // @[LZD.scala 39:27]
  assign _T_79 = _T_76 | _T_78; // @[LZD.scala 39:25]
  assign _T_80 = {_T_75,_T_79}; // @[Cat.scala 29:58]
  assign _T_81 = _T_73[1:0]; // @[LZD.scala 44:32]
  assign _T_82 = _T_81 != 2'h0; // @[LZD.scala 39:14]
  assign _T_83 = _T_81[1]; // @[LZD.scala 39:21]
  assign _T_84 = _T_81[0]; // @[LZD.scala 39:30]
  assign _T_85 = ~ _T_84; // @[LZD.scala 39:27]
  assign _T_86 = _T_83 | _T_85; // @[LZD.scala 39:25]
  assign _T_87 = {_T_82,_T_86}; // @[Cat.scala 29:58]
  assign _T_88 = _T_80[1]; // @[Shift.scala 12:21]
  assign _T_89 = _T_87[1]; // @[Shift.scala 12:21]
  assign _T_90 = _T_88 | _T_89; // @[LZD.scala 49:16]
  assign _T_91 = ~ _T_89; // @[LZD.scala 49:27]
  assign _T_92 = _T_88 | _T_91; // @[LZD.scala 49:25]
  assign _T_93 = _T_80[0:0]; // @[LZD.scala 49:47]
  assign _T_94 = _T_87[0:0]; // @[LZD.scala 49:59]
  assign _T_95 = _T_88 ? _T_93 : _T_94; // @[LZD.scala 49:35]
  assign _T_97 = {_T_90,_T_92,_T_95}; // @[Cat.scala 29:58]
  assign _T_98 = _T_72[3:0]; // @[LZD.scala 44:32]
  assign _T_99 = _T_98[3:2]; // @[LZD.scala 43:32]
  assign _T_100 = _T_99 != 2'h0; // @[LZD.scala 39:14]
  assign _T_101 = _T_99[1]; // @[LZD.scala 39:21]
  assign _T_102 = _T_99[0]; // @[LZD.scala 39:30]
  assign _T_103 = ~ _T_102; // @[LZD.scala 39:27]
  assign _T_104 = _T_101 | _T_103; // @[LZD.scala 39:25]
  assign _T_105 = {_T_100,_T_104}; // @[Cat.scala 29:58]
  assign _T_106 = _T_98[1:0]; // @[LZD.scala 44:32]
  assign _T_107 = _T_106 != 2'h0; // @[LZD.scala 39:14]
  assign _T_108 = _T_106[1]; // @[LZD.scala 39:21]
  assign _T_109 = _T_106[0]; // @[LZD.scala 39:30]
  assign _T_110 = ~ _T_109; // @[LZD.scala 39:27]
  assign _T_111 = _T_108 | _T_110; // @[LZD.scala 39:25]
  assign _T_112 = {_T_107,_T_111}; // @[Cat.scala 29:58]
  assign _T_113 = _T_105[1]; // @[Shift.scala 12:21]
  assign _T_114 = _T_112[1]; // @[Shift.scala 12:21]
  assign _T_115 = _T_113 | _T_114; // @[LZD.scala 49:16]
  assign _T_116 = ~ _T_114; // @[LZD.scala 49:27]
  assign _T_117 = _T_113 | _T_116; // @[LZD.scala 49:25]
  assign _T_118 = _T_105[0:0]; // @[LZD.scala 49:47]
  assign _T_119 = _T_112[0:0]; // @[LZD.scala 49:59]
  assign _T_120 = _T_113 ? _T_118 : _T_119; // @[LZD.scala 49:35]
  assign _T_122 = {_T_115,_T_117,_T_120}; // @[Cat.scala 29:58]
  assign _T_123 = _T_97[2]; // @[Shift.scala 12:21]
  assign _T_124 = _T_122[2]; // @[Shift.scala 12:21]
  assign _T_125 = _T_123 | _T_124; // @[LZD.scala 49:16]
  assign _T_126 = ~ _T_124; // @[LZD.scala 49:27]
  assign _T_127 = _T_123 | _T_126; // @[LZD.scala 49:25]
  assign _T_128 = _T_97[1:0]; // @[LZD.scala 49:47]
  assign _T_129 = _T_122[1:0]; // @[LZD.scala 49:59]
  assign _T_130 = _T_123 ? _T_128 : _T_129; // @[LZD.scala 49:35]
  assign _T_132 = {_T_125,_T_127,_T_130}; // @[Cat.scala 29:58]
  assign _T_133 = _T_71[3]; // @[Shift.scala 12:21]
  assign _T_134 = _T_132[3]; // @[Shift.scala 12:21]
  assign _T_135 = _T_133 | _T_134; // @[LZD.scala 49:16]
  assign _T_136 = ~ _T_134; // @[LZD.scala 49:27]
  assign _T_137 = _T_133 | _T_136; // @[LZD.scala 49:25]
  assign _T_138 = _T_71[2:0]; // @[LZD.scala 49:47]
  assign _T_139 = _T_132[2:0]; // @[LZD.scala 49:59]
  assign _T_140 = _T_133 ? _T_138 : _T_139; // @[LZD.scala 49:35]
  assign _T_142 = {_T_135,_T_137,_T_140}; // @[Cat.scala 29:58]
  assign _T_143 = quireXOR[14:0]; // @[LZD.scala 44:32]
  assign _T_144 = _T_143[14:7]; // @[LZD.scala 43:32]
  assign _T_145 = _T_144[7:4]; // @[LZD.scala 43:32]
  assign _T_146 = _T_145[3:2]; // @[LZD.scala 43:32]
  assign _T_147 = _T_146 != 2'h0; // @[LZD.scala 39:14]
  assign _T_148 = _T_146[1]; // @[LZD.scala 39:21]
  assign _T_149 = _T_146[0]; // @[LZD.scala 39:30]
  assign _T_150 = ~ _T_149; // @[LZD.scala 39:27]
  assign _T_151 = _T_148 | _T_150; // @[LZD.scala 39:25]
  assign _T_152 = {_T_147,_T_151}; // @[Cat.scala 29:58]
  assign _T_153 = _T_145[1:0]; // @[LZD.scala 44:32]
  assign _T_154 = _T_153 != 2'h0; // @[LZD.scala 39:14]
  assign _T_155 = _T_153[1]; // @[LZD.scala 39:21]
  assign _T_156 = _T_153[0]; // @[LZD.scala 39:30]
  assign _T_157 = ~ _T_156; // @[LZD.scala 39:27]
  assign _T_158 = _T_155 | _T_157; // @[LZD.scala 39:25]
  assign _T_159 = {_T_154,_T_158}; // @[Cat.scala 29:58]
  assign _T_160 = _T_152[1]; // @[Shift.scala 12:21]
  assign _T_161 = _T_159[1]; // @[Shift.scala 12:21]
  assign _T_162 = _T_160 | _T_161; // @[LZD.scala 49:16]
  assign _T_163 = ~ _T_161; // @[LZD.scala 49:27]
  assign _T_164 = _T_160 | _T_163; // @[LZD.scala 49:25]
  assign _T_165 = _T_152[0:0]; // @[LZD.scala 49:47]
  assign _T_166 = _T_159[0:0]; // @[LZD.scala 49:59]
  assign _T_167 = _T_160 ? _T_165 : _T_166; // @[LZD.scala 49:35]
  assign _T_169 = {_T_162,_T_164,_T_167}; // @[Cat.scala 29:58]
  assign _T_170 = _T_144[3:0]; // @[LZD.scala 44:32]
  assign _T_171 = _T_170[3:2]; // @[LZD.scala 43:32]
  assign _T_172 = _T_171 != 2'h0; // @[LZD.scala 39:14]
  assign _T_173 = _T_171[1]; // @[LZD.scala 39:21]
  assign _T_174 = _T_171[0]; // @[LZD.scala 39:30]
  assign _T_175 = ~ _T_174; // @[LZD.scala 39:27]
  assign _T_176 = _T_173 | _T_175; // @[LZD.scala 39:25]
  assign _T_177 = {_T_172,_T_176}; // @[Cat.scala 29:58]
  assign _T_178 = _T_170[1:0]; // @[LZD.scala 44:32]
  assign _T_179 = _T_178 != 2'h0; // @[LZD.scala 39:14]
  assign _T_180 = _T_178[1]; // @[LZD.scala 39:21]
  assign _T_181 = _T_178[0]; // @[LZD.scala 39:30]
  assign _T_182 = ~ _T_181; // @[LZD.scala 39:27]
  assign _T_183 = _T_180 | _T_182; // @[LZD.scala 39:25]
  assign _T_184 = {_T_179,_T_183}; // @[Cat.scala 29:58]
  assign _T_185 = _T_177[1]; // @[Shift.scala 12:21]
  assign _T_186 = _T_184[1]; // @[Shift.scala 12:21]
  assign _T_187 = _T_185 | _T_186; // @[LZD.scala 49:16]
  assign _T_188 = ~ _T_186; // @[LZD.scala 49:27]
  assign _T_189 = _T_185 | _T_188; // @[LZD.scala 49:25]
  assign _T_190 = _T_177[0:0]; // @[LZD.scala 49:47]
  assign _T_191 = _T_184[0:0]; // @[LZD.scala 49:59]
  assign _T_192 = _T_185 ? _T_190 : _T_191; // @[LZD.scala 49:35]
  assign _T_194 = {_T_187,_T_189,_T_192}; // @[Cat.scala 29:58]
  assign _T_195 = _T_169[2]; // @[Shift.scala 12:21]
  assign _T_196 = _T_194[2]; // @[Shift.scala 12:21]
  assign _T_197 = _T_195 | _T_196; // @[LZD.scala 49:16]
  assign _T_198 = ~ _T_196; // @[LZD.scala 49:27]
  assign _T_199 = _T_195 | _T_198; // @[LZD.scala 49:25]
  assign _T_200 = _T_169[1:0]; // @[LZD.scala 49:47]
  assign _T_201 = _T_194[1:0]; // @[LZD.scala 49:59]
  assign _T_202 = _T_195 ? _T_200 : _T_201; // @[LZD.scala 49:35]
  assign _T_204 = {_T_197,_T_199,_T_202}; // @[Cat.scala 29:58]
  assign _T_205 = _T_143[6:0]; // @[LZD.scala 44:32]
  assign _T_206 = _T_205[6:3]; // @[LZD.scala 43:32]
  assign _T_207 = _T_206[3:2]; // @[LZD.scala 43:32]
  assign _T_208 = _T_207 != 2'h0; // @[LZD.scala 39:14]
  assign _T_209 = _T_207[1]; // @[LZD.scala 39:21]
  assign _T_210 = _T_207[0]; // @[LZD.scala 39:30]
  assign _T_211 = ~ _T_210; // @[LZD.scala 39:27]
  assign _T_212 = _T_209 | _T_211; // @[LZD.scala 39:25]
  assign _T_213 = {_T_208,_T_212}; // @[Cat.scala 29:58]
  assign _T_214 = _T_206[1:0]; // @[LZD.scala 44:32]
  assign _T_215 = _T_214 != 2'h0; // @[LZD.scala 39:14]
  assign _T_216 = _T_214[1]; // @[LZD.scala 39:21]
  assign _T_217 = _T_214[0]; // @[LZD.scala 39:30]
  assign _T_218 = ~ _T_217; // @[LZD.scala 39:27]
  assign _T_219 = _T_216 | _T_218; // @[LZD.scala 39:25]
  assign _T_220 = {_T_215,_T_219}; // @[Cat.scala 29:58]
  assign _T_221 = _T_213[1]; // @[Shift.scala 12:21]
  assign _T_222 = _T_220[1]; // @[Shift.scala 12:21]
  assign _T_223 = _T_221 | _T_222; // @[LZD.scala 49:16]
  assign _T_224 = ~ _T_222; // @[LZD.scala 49:27]
  assign _T_225 = _T_221 | _T_224; // @[LZD.scala 49:25]
  assign _T_226 = _T_213[0:0]; // @[LZD.scala 49:47]
  assign _T_227 = _T_220[0:0]; // @[LZD.scala 49:59]
  assign _T_228 = _T_221 ? _T_226 : _T_227; // @[LZD.scala 49:35]
  assign _T_230 = {_T_223,_T_225,_T_228}; // @[Cat.scala 29:58]
  assign _T_231 = _T_205[2:0]; // @[LZD.scala 44:32]
  assign _T_232 = _T_231[2:1]; // @[LZD.scala 43:32]
  assign _T_233 = _T_232 != 2'h0; // @[LZD.scala 39:14]
  assign _T_234 = _T_232[1]; // @[LZD.scala 39:21]
  assign _T_235 = _T_232[0]; // @[LZD.scala 39:30]
  assign _T_236 = ~ _T_235; // @[LZD.scala 39:27]
  assign _T_237 = _T_234 | _T_236; // @[LZD.scala 39:25]
  assign _T_238 = {_T_233,_T_237}; // @[Cat.scala 29:58]
  assign _T_239 = _T_231[0:0]; // @[LZD.scala 44:32]
  assign _T_241 = _T_238[1]; // @[Shift.scala 12:21]
  assign _T_243 = _T_238[0:0]; // @[LZD.scala 55:32]
  assign _T_244 = _T_241 ? _T_243 : _T_239; // @[LZD.scala 55:20]
  assign _T_245 = {_T_241,_T_244}; // @[Cat.scala 29:58]
  assign _T_246 = _T_230[2]; // @[Shift.scala 12:21]
  assign _T_248 = _T_230[1:0]; // @[LZD.scala 55:32]
  assign _T_249 = _T_246 ? _T_248 : _T_245; // @[LZD.scala 55:20]
  assign _T_250 = {_T_246,_T_249}; // @[Cat.scala 29:58]
  assign _T_251 = _T_204[3]; // @[Shift.scala 12:21]
  assign _T_253 = _T_204[2:0]; // @[LZD.scala 55:32]
  assign _T_254 = _T_251 ? _T_253 : _T_250; // @[LZD.scala 55:20]
  assign _T_255 = {_T_251,_T_254}; // @[Cat.scala 29:58]
  assign _T_256 = _T_142[4]; // @[Shift.scala 12:21]
  assign _T_258 = _T_142[3:0]; // @[LZD.scala 55:32]
  assign _T_259 = _T_256 ? _T_258 : _T_255; // @[LZD.scala 55:20]
  assign scaleBias = {1'h1,_T_256,_T_259}; // @[Cat.scala 29:58]
  assign _T_260 = $signed(scaleBias); // @[QuireToPosit.scala 61:53]
  assign _GEN_2 = {{1{_T_260[5]}},_T_260}; // @[QuireToPosit.scala 61:41]
  assign _T_262 = $signed(7'sh13) + $signed(_GEN_2); // @[QuireToPosit.scala 61:41]
  assign realScale = $signed(_T_262); // @[QuireToPosit.scala 61:41]
  assign underflow = $signed(realScale) < $signed(-7'sh7); // @[QuireToPosit.scala 62:41]
  assign overflow = $signed(realScale) > $signed(7'sh6); // @[QuireToPosit.scala 63:35]
  assign _T_263 = underflow ? $signed(-7'sh7) : $signed(realScale); // @[Mux.scala 87:16]
  assign _T_264 = overflow ? $signed(7'sh6) : $signed(_T_263); // @[Mux.scala 87:16]
  assign _T_265 = realScale[6:6]; // @[Abs.scala 10:21]
  assign _T_267 = _T_265 ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign _T_268 = $unsigned(realScale); // @[Abs.scala 10:31]
  assign _T_269 = _T_267 ^ _T_268; // @[Abs.scala 10:26]
  assign _GEN_3 = {{6'd0}, _T_265}; // @[Abs.scala 10:39]
  assign absRealScale = _T_269 + _GEN_3; // @[Abs.scala 10:39]
  assign _T_272 = absRealScale < 7'h20; // @[Shift.scala 16:24]
  assign _T_273 = absRealScale[4:0]; // @[Shift.scala 17:37]
  assign _T_274 = _T_273[4]; // @[Shift.scala 12:21]
  assign _T_275 = io_quireIn[15:0]; // @[Shift.scala 64:52]
  assign _T_277 = {_T_275,16'h0}; // @[Cat.scala 29:58]
  assign _T_278 = _T_274 ? _T_277 : io_quireIn; // @[Shift.scala 64:27]
  assign _T_279 = _T_273[3:0]; // @[Shift.scala 66:70]
  assign _T_280 = _T_279[3]; // @[Shift.scala 12:21]
  assign _T_281 = _T_278[23:0]; // @[Shift.scala 64:52]
  assign _T_283 = {_T_281,8'h0}; // @[Cat.scala 29:58]
  assign _T_284 = _T_280 ? _T_283 : _T_278; // @[Shift.scala 64:27]
  assign _T_285 = _T_279[2:0]; // @[Shift.scala 66:70]
  assign _T_286 = _T_285[2]; // @[Shift.scala 12:21]
  assign _T_287 = _T_284[27:0]; // @[Shift.scala 64:52]
  assign _T_289 = {_T_287,4'h0}; // @[Cat.scala 29:58]
  assign _T_290 = _T_286 ? _T_289 : _T_284; // @[Shift.scala 64:27]
  assign _T_291 = _T_285[1:0]; // @[Shift.scala 66:70]
  assign _T_292 = _T_291[1]; // @[Shift.scala 12:21]
  assign _T_293 = _T_290[29:0]; // @[Shift.scala 64:52]
  assign _T_295 = {_T_293,2'h0}; // @[Cat.scala 29:58]
  assign _T_296 = _T_292 ? _T_295 : _T_290; // @[Shift.scala 64:27]
  assign _T_297 = _T_291[0:0]; // @[Shift.scala 66:70]
  assign _T_299 = _T_296[30:0]; // @[Shift.scala 64:52]
  assign _T_300 = {_T_299,1'h0}; // @[Cat.scala 29:58]
  assign _T_301 = _T_297 ? _T_300 : _T_296; // @[Shift.scala 64:27]
  assign quireLeftShift = _T_272 ? _T_301 : 32'h0; // @[Shift.scala 16:10]
  assign _T_306 = io_quireIn[31:16]; // @[Shift.scala 77:66]
  assign _T_307 = {16'h0,_T_306}; // @[Cat.scala 29:58]
  assign _T_308 = _T_274 ? _T_307 : io_quireIn; // @[Shift.scala 77:22]
  assign _T_312 = _T_308[31:8]; // @[Shift.scala 77:66]
  assign _T_313 = {8'h0,_T_312}; // @[Cat.scala 29:58]
  assign _T_314 = _T_280 ? _T_313 : _T_308; // @[Shift.scala 77:22]
  assign _T_318 = _T_314[31:4]; // @[Shift.scala 77:66]
  assign _T_319 = {4'h0,_T_318}; // @[Cat.scala 29:58]
  assign _T_320 = _T_286 ? _T_319 : _T_314; // @[Shift.scala 77:22]
  assign _T_324 = _T_320[31:2]; // @[Shift.scala 77:66]
  assign _T_325 = {2'h0,_T_324}; // @[Cat.scala 29:58]
  assign _T_326 = _T_292 ? _T_325 : _T_320; // @[Shift.scala 77:22]
  assign _T_329 = _T_326[31:1]; // @[Shift.scala 77:66]
  assign _T_330 = {1'h0,_T_329}; // @[Cat.scala 29:58]
  assign _T_331 = _T_297 ? _T_330 : _T_326; // @[Shift.scala 77:22]
  assign quireRightShift = _T_272 ? _T_331 : 32'h0; // @[Shift.scala 27:10]
  assign _T_333 = quireLeftShift[11:5]; // @[QuireToPosit.scala 89:49]
  assign _T_334 = quireLeftShift[4:0]; // @[QuireToPosit.scala 90:127]
  assign _T_335 = _T_334 != 5'h0; // @[QuireToPosit.scala 90:154]
  assign realFGRSTmp1 = {_T_333,_T_335}; // @[Cat.scala 29:58]
  assign _T_336 = quireRightShift[11:5]; // @[QuireToPosit.scala 91:50]
  assign _T_337 = quireRightShift[4:0]; // @[QuireToPosit.scala 92:128]
  assign _T_338 = _T_337 != 5'h0; // @[QuireToPosit.scala 92:155]
  assign realFGRSTmp2 = {_T_336,_T_338}; // @[Cat.scala 29:58]
  assign realFGRS = _T_265 ? realFGRSTmp1 : realFGRSTmp2; // @[QuireToPosit.scala 93:34]
  assign outRawFloat_fraction = realFGRS[7:3]; // @[QuireToPosit.scala 95:46]
  assign outRawFloat_grs = realFGRS[2:0]; // @[QuireToPosit.scala 96:46]
  assign _GEN_4 = _T_264[3:0]; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  assign outRawFloat_scale = $signed(_GEN_4); // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  assign _T_344 = outRawFloat_scale[3:3]; // @[convert.scala 49:36]
  assign _T_346 = ~ outRawFloat_scale; // @[convert.scala 50:36]
  assign _T_347 = $signed(_T_346); // @[convert.scala 50:36]
  assign _T_348 = _T_344 ? $signed(_T_347) : $signed(outRawFloat_scale); // @[convert.scala 50:28]
  assign _T_349 = _T_344 ^ _T_2; // @[convert.scala 51:31]
  assign _T_350 = ~ _T_349; // @[convert.scala 53:34]
  assign _T_353 = {_T_350,_T_349,outRawFloat_fraction,outRawFloat_grs}; // @[Cat.scala 29:58]
  assign _T_354 = $unsigned(_T_348); // @[Shift.scala 39:17]
  assign _T_355 = _T_354 < 4'ha; // @[Shift.scala 39:24]
  assign _T_357 = _T_353[9:8]; // @[Shift.scala 90:30]
  assign _T_358 = _T_353[7:0]; // @[Shift.scala 90:48]
  assign _T_359 = _T_358 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{1'd0}, _T_359}; // @[Shift.scala 90:39]
  assign _T_360 = _T_357 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_361 = _T_354[3]; // @[Shift.scala 12:21]
  assign _T_362 = _T_353[9]; // @[Shift.scala 12:21]
  assign _T_364 = _T_362 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_365 = {_T_364,_T_360}; // @[Cat.scala 29:58]
  assign _T_366 = _T_361 ? _T_365 : _T_353; // @[Shift.scala 91:22]
  assign _T_367 = _T_354[2:0]; // @[Shift.scala 92:77]
  assign _T_368 = _T_366[9:4]; // @[Shift.scala 90:30]
  assign _T_369 = _T_366[3:0]; // @[Shift.scala 90:48]
  assign _T_370 = _T_369 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{5'd0}, _T_370}; // @[Shift.scala 90:39]
  assign _T_371 = _T_368 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_372 = _T_367[2]; // @[Shift.scala 12:21]
  assign _T_373 = _T_366[9]; // @[Shift.scala 12:21]
  assign _T_375 = _T_373 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_376 = {_T_375,_T_371}; // @[Cat.scala 29:58]
  assign _T_377 = _T_372 ? _T_376 : _T_366; // @[Shift.scala 91:22]
  assign _T_378 = _T_367[1:0]; // @[Shift.scala 92:77]
  assign _T_379 = _T_377[9:2]; // @[Shift.scala 90:30]
  assign _T_380 = _T_377[1:0]; // @[Shift.scala 90:48]
  assign _T_381 = _T_380 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{7'd0}, _T_381}; // @[Shift.scala 90:39]
  assign _T_382 = _T_379 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_383 = _T_378[1]; // @[Shift.scala 12:21]
  assign _T_384 = _T_377[9]; // @[Shift.scala 12:21]
  assign _T_386 = _T_384 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_387 = {_T_386,_T_382}; // @[Cat.scala 29:58]
  assign _T_388 = _T_383 ? _T_387 : _T_377; // @[Shift.scala 91:22]
  assign _T_389 = _T_378[0:0]; // @[Shift.scala 92:77]
  assign _T_390 = _T_388[9:1]; // @[Shift.scala 90:30]
  assign _T_391 = _T_388[0:0]; // @[Shift.scala 90:48]
  assign _GEN_8 = {{8'd0}, _T_391}; // @[Shift.scala 90:39]
  assign _T_393 = _T_390 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_395 = _T_388[9]; // @[Shift.scala 12:21]
  assign _T_396 = {_T_395,_T_393}; // @[Cat.scala 29:58]
  assign _T_397 = _T_389 ? _T_396 : _T_388; // @[Shift.scala 91:22]
  assign _T_400 = _T_362 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_401 = _T_355 ? _T_397 : _T_400; // @[Shift.scala 39:10]
  assign _T_402 = _T_401[3]; // @[convert.scala 55:31]
  assign _T_403 = _T_401[2]; // @[convert.scala 56:31]
  assign _T_404 = _T_401[1]; // @[convert.scala 57:31]
  assign _T_405 = _T_401[0]; // @[convert.scala 58:31]
  assign _T_406 = _T_401[9:3]; // @[convert.scala 59:69]
  assign _T_407 = _T_406 != 7'h0; // @[convert.scala 59:81]
  assign _T_408 = ~ _T_407; // @[convert.scala 59:50]
  assign _T_410 = _T_406 == 7'h7f; // @[convert.scala 60:81]
  assign _T_411 = _T_402 | _T_404; // @[convert.scala 61:44]
  assign _T_412 = _T_411 | _T_405; // @[convert.scala 61:52]
  assign _T_413 = _T_403 & _T_412; // @[convert.scala 61:36]
  assign _T_414 = ~ _T_410; // @[convert.scala 62:63]
  assign _T_415 = _T_414 & _T_413; // @[convert.scala 62:103]
  assign _T_416 = _T_408 | _T_415; // @[convert.scala 62:60]
  assign _GEN_9 = {{6'd0}, _T_416}; // @[convert.scala 63:56]
  assign _T_419 = _T_406 + _GEN_9; // @[convert.scala 63:56]
  assign _T_420 = {_T_2,_T_419}; // @[Cat.scala 29:58]
  assign io_positOut = _T_428; // @[QuireToPosit.scala 101:15]
  assign io_outValid = _T_424; // @[QuireToPosit.scala 100:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_424 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_428 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_424 <= 1'h0;
    end else begin
      _T_424 <= io_inValid;
    end
    if (io_inValid) begin
      if (outRawFloat_isNaR) begin
        _T_428 <= 8'h80;
      end else begin
        if (outRawFloat_isZero) begin
          _T_428 <= 8'h0;
        end else begin
          _T_428 <= _T_420;
        end
      end
    end
  end
endmodule
