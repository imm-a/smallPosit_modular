module QuireToPosit6_4_0(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [15:0] io_quireIn,
  output [3:0]  io_positOut,
  output        io_outValid
);
  wire [14:0] _T; // @[QuireToPosit.scala 47:43]
  wire  _T_1; // @[QuireToPosit.scala 47:47]
  wire  tailIsZero; // @[QuireToPosit.scala 47:27]
  wire  _T_2; // @[QuireToPosit.scala 49:45]
  wire  outRawFloat_isNaR; // @[QuireToPosit.scala 49:49]
  wire  _T_5; // @[QuireToPosit.scala 50:31]
  wire  outRawFloat_isZero; // @[QuireToPosit.scala 50:51]
  wire [14:0] _T_8; // @[QuireToPosit.scala 58:41]
  wire [14:0] _T_9; // @[QuireToPosit.scala 58:68]
  wire [14:0] quireXOR; // @[QuireToPosit.scala 58:56]
  wire [7:0] _T_10; // @[LZD.scala 43:32]
  wire [3:0] _T_11; // @[LZD.scala 43:32]
  wire [1:0] _T_12; // @[LZD.scala 43:32]
  wire  _T_13; // @[LZD.scala 39:14]
  wire  _T_14; // @[LZD.scala 39:21]
  wire  _T_15; // @[LZD.scala 39:30]
  wire  _T_16; // @[LZD.scala 39:27]
  wire  _T_17; // @[LZD.scala 39:25]
  wire [1:0] _T_18; // @[Cat.scala 29:58]
  wire [1:0] _T_19; // @[LZD.scala 44:32]
  wire  _T_20; // @[LZD.scala 39:14]
  wire  _T_21; // @[LZD.scala 39:21]
  wire  _T_22; // @[LZD.scala 39:30]
  wire  _T_23; // @[LZD.scala 39:27]
  wire  _T_24; // @[LZD.scala 39:25]
  wire [1:0] _T_25; // @[Cat.scala 29:58]
  wire  _T_26; // @[Shift.scala 12:21]
  wire  _T_27; // @[Shift.scala 12:21]
  wire  _T_28; // @[LZD.scala 49:16]
  wire  _T_29; // @[LZD.scala 49:27]
  wire  _T_30; // @[LZD.scala 49:25]
  wire  _T_31; // @[LZD.scala 49:47]
  wire  _T_32; // @[LZD.scala 49:59]
  wire  _T_33; // @[LZD.scala 49:35]
  wire [2:0] _T_35; // @[Cat.scala 29:58]
  wire [3:0] _T_36; // @[LZD.scala 44:32]
  wire [1:0] _T_37; // @[LZD.scala 43:32]
  wire  _T_38; // @[LZD.scala 39:14]
  wire  _T_39; // @[LZD.scala 39:21]
  wire  _T_40; // @[LZD.scala 39:30]
  wire  _T_41; // @[LZD.scala 39:27]
  wire  _T_42; // @[LZD.scala 39:25]
  wire [1:0] _T_43; // @[Cat.scala 29:58]
  wire [1:0] _T_44; // @[LZD.scala 44:32]
  wire  _T_45; // @[LZD.scala 39:14]
  wire  _T_46; // @[LZD.scala 39:21]
  wire  _T_47; // @[LZD.scala 39:30]
  wire  _T_48; // @[LZD.scala 39:27]
  wire  _T_49; // @[LZD.scala 39:25]
  wire [1:0] _T_50; // @[Cat.scala 29:58]
  wire  _T_51; // @[Shift.scala 12:21]
  wire  _T_52; // @[Shift.scala 12:21]
  wire  _T_53; // @[LZD.scala 49:16]
  wire  _T_54; // @[LZD.scala 49:27]
  wire  _T_55; // @[LZD.scala 49:25]
  wire  _T_56; // @[LZD.scala 49:47]
  wire  _T_57; // @[LZD.scala 49:59]
  wire  _T_58; // @[LZD.scala 49:35]
  wire [2:0] _T_60; // @[Cat.scala 29:58]
  wire  _T_61; // @[Shift.scala 12:21]
  wire  _T_62; // @[Shift.scala 12:21]
  wire  _T_63; // @[LZD.scala 49:16]
  wire  _T_64; // @[LZD.scala 49:27]
  wire  _T_65; // @[LZD.scala 49:25]
  wire [1:0] _T_66; // @[LZD.scala 49:47]
  wire [1:0] _T_67; // @[LZD.scala 49:59]
  wire [1:0] _T_68; // @[LZD.scala 49:35]
  wire [3:0] _T_70; // @[Cat.scala 29:58]
  wire [6:0] _T_71; // @[LZD.scala 44:32]
  wire [3:0] _T_72; // @[LZD.scala 43:32]
  wire [1:0] _T_73; // @[LZD.scala 43:32]
  wire  _T_74; // @[LZD.scala 39:14]
  wire  _T_75; // @[LZD.scala 39:21]
  wire  _T_76; // @[LZD.scala 39:30]
  wire  _T_77; // @[LZD.scala 39:27]
  wire  _T_78; // @[LZD.scala 39:25]
  wire [1:0] _T_79; // @[Cat.scala 29:58]
  wire [1:0] _T_80; // @[LZD.scala 44:32]
  wire  _T_81; // @[LZD.scala 39:14]
  wire  _T_82; // @[LZD.scala 39:21]
  wire  _T_83; // @[LZD.scala 39:30]
  wire  _T_84; // @[LZD.scala 39:27]
  wire  _T_85; // @[LZD.scala 39:25]
  wire [1:0] _T_86; // @[Cat.scala 29:58]
  wire  _T_87; // @[Shift.scala 12:21]
  wire  _T_88; // @[Shift.scala 12:21]
  wire  _T_89; // @[LZD.scala 49:16]
  wire  _T_90; // @[LZD.scala 49:27]
  wire  _T_91; // @[LZD.scala 49:25]
  wire  _T_92; // @[LZD.scala 49:47]
  wire  _T_93; // @[LZD.scala 49:59]
  wire  _T_94; // @[LZD.scala 49:35]
  wire [2:0] _T_96; // @[Cat.scala 29:58]
  wire [2:0] _T_97; // @[LZD.scala 44:32]
  wire [1:0] _T_98; // @[LZD.scala 43:32]
  wire  _T_99; // @[LZD.scala 39:14]
  wire  _T_100; // @[LZD.scala 39:21]
  wire  _T_101; // @[LZD.scala 39:30]
  wire  _T_102; // @[LZD.scala 39:27]
  wire  _T_103; // @[LZD.scala 39:25]
  wire [1:0] _T_104; // @[Cat.scala 29:58]
  wire  _T_105; // @[LZD.scala 44:32]
  wire  _T_107; // @[Shift.scala 12:21]
  wire  _T_109; // @[LZD.scala 55:32]
  wire  _T_110; // @[LZD.scala 55:20]
  wire [1:0] _T_111; // @[Cat.scala 29:58]
  wire  _T_112; // @[Shift.scala 12:21]
  wire [1:0] _T_114; // @[LZD.scala 55:32]
  wire [1:0] _T_115; // @[LZD.scala 55:20]
  wire [2:0] _T_116; // @[Cat.scala 29:58]
  wire  _T_117; // @[Shift.scala 12:21]
  wire [2:0] _T_119; // @[LZD.scala 55:32]
  wire [2:0] _T_120; // @[LZD.scala 55:20]
  wire [4:0] scaleBias; // @[Cat.scala 29:58]
  wire [4:0] _T_121; // @[QuireToPosit.scala 61:53]
  wire [5:0] _GEN_2; // @[QuireToPosit.scala 61:41]
  wire [5:0] _T_123; // @[QuireToPosit.scala 61:41]
  wire [5:0] realScale; // @[QuireToPosit.scala 61:41]
  wire  underflow; // @[QuireToPosit.scala 62:41]
  wire  overflow; // @[QuireToPosit.scala 63:35]
  wire [5:0] _T_124; // @[Mux.scala 87:16]
  wire [5:0] _T_125; // @[Mux.scala 87:16]
  wire  _T_126; // @[Abs.scala 10:21]
  wire [5:0] _T_128; // @[Bitwise.scala 71:12]
  wire [5:0] _T_129; // @[Abs.scala 10:31]
  wire [5:0] _T_130; // @[Abs.scala 10:26]
  wire [5:0] _GEN_3; // @[Abs.scala 10:39]
  wire [5:0] absRealScale; // @[Abs.scala 10:39]
  wire  _T_133; // @[Shift.scala 16:24]
  wire [3:0] _T_134; // @[Shift.scala 17:37]
  wire  _T_135; // @[Shift.scala 12:21]
  wire [7:0] _T_136; // @[Shift.scala 64:52]
  wire [15:0] _T_138; // @[Cat.scala 29:58]
  wire [15:0] _T_139; // @[Shift.scala 64:27]
  wire [2:0] _T_140; // @[Shift.scala 66:70]
  wire  _T_141; // @[Shift.scala 12:21]
  wire [11:0] _T_142; // @[Shift.scala 64:52]
  wire [15:0] _T_144; // @[Cat.scala 29:58]
  wire [15:0] _T_145; // @[Shift.scala 64:27]
  wire [1:0] _T_146; // @[Shift.scala 66:70]
  wire  _T_147; // @[Shift.scala 12:21]
  wire [13:0] _T_148; // @[Shift.scala 64:52]
  wire [15:0] _T_150; // @[Cat.scala 29:58]
  wire [15:0] _T_151; // @[Shift.scala 64:27]
  wire  _T_152; // @[Shift.scala 66:70]
  wire [14:0] _T_154; // @[Shift.scala 64:52]
  wire [15:0] _T_155; // @[Cat.scala 29:58]
  wire [15:0] _T_156; // @[Shift.scala 64:27]
  wire [15:0] quireLeftShift; // @[Shift.scala 16:10]
  wire [7:0] _T_161; // @[Shift.scala 77:66]
  wire [15:0] _T_162; // @[Cat.scala 29:58]
  wire [15:0] _T_163; // @[Shift.scala 77:22]
  wire [11:0] _T_167; // @[Shift.scala 77:66]
  wire [15:0] _T_168; // @[Cat.scala 29:58]
  wire [15:0] _T_169; // @[Shift.scala 77:22]
  wire [13:0] _T_173; // @[Shift.scala 77:66]
  wire [15:0] _T_174; // @[Cat.scala 29:58]
  wire [15:0] _T_175; // @[Shift.scala 77:22]
  wire [14:0] _T_178; // @[Shift.scala 77:66]
  wire [15:0] _T_179; // @[Cat.scala 29:58]
  wire [15:0] _T_180; // @[Shift.scala 77:22]
  wire [15:0] quireRightShift; // @[Shift.scala 27:10]
  wire [2:0] _T_182; // @[QuireToPosit.scala 89:49]
  wire  _T_183; // @[QuireToPosit.scala 90:127]
  wire [3:0] realFGRSTmp1; // @[Cat.scala 29:58]
  wire [2:0] _T_185; // @[QuireToPosit.scala 91:50]
  wire  _T_186; // @[QuireToPosit.scala 92:128]
  wire [3:0] realFGRSTmp2; // @[Cat.scala 29:58]
  wire [3:0] realFGRS; // @[QuireToPosit.scala 93:34]
  wire  outRawFloat_fraction; // @[QuireToPosit.scala 95:46]
  wire [2:0] outRawFloat_grs; // @[QuireToPosit.scala 96:46]
  wire [2:0] _GEN_4; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  wire [2:0] outRawFloat_scale; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  wire  _T_193; // @[convert.scala 49:36]
  wire [2:0] _T_195; // @[convert.scala 50:36]
  wire [2:0] _T_196; // @[convert.scala 50:36]
  wire [2:0] _T_197; // @[convert.scala 50:28]
  wire  _T_198; // @[convert.scala 51:31]
  wire  _T_199; // @[convert.scala 53:34]
  wire [5:0] _T_202; // @[Cat.scala 29:58]
  wire [2:0] _T_203; // @[Shift.scala 39:17]
  wire  _T_204; // @[Shift.scala 39:24]
  wire [1:0] _T_206; // @[Shift.scala 90:30]
  wire [3:0] _T_207; // @[Shift.scala 90:48]
  wire  _T_208; // @[Shift.scala 90:57]
  wire [1:0] _GEN_5; // @[Shift.scala 90:39]
  wire [1:0] _T_209; // @[Shift.scala 90:39]
  wire  _T_210; // @[Shift.scala 12:21]
  wire  _T_211; // @[Shift.scala 12:21]
  wire [3:0] _T_213; // @[Bitwise.scala 71:12]
  wire [5:0] _T_214; // @[Cat.scala 29:58]
  wire [5:0] _T_215; // @[Shift.scala 91:22]
  wire [1:0] _T_216; // @[Shift.scala 92:77]
  wire [3:0] _T_217; // @[Shift.scala 90:30]
  wire [1:0] _T_218; // @[Shift.scala 90:48]
  wire  _T_219; // @[Shift.scala 90:57]
  wire [3:0] _GEN_6; // @[Shift.scala 90:39]
  wire [3:0] _T_220; // @[Shift.scala 90:39]
  wire  _T_221; // @[Shift.scala 12:21]
  wire  _T_222; // @[Shift.scala 12:21]
  wire [1:0] _T_224; // @[Bitwise.scala 71:12]
  wire [5:0] _T_225; // @[Cat.scala 29:58]
  wire [5:0] _T_226; // @[Shift.scala 91:22]
  wire  _T_227; // @[Shift.scala 92:77]
  wire [4:0] _T_228; // @[Shift.scala 90:30]
  wire  _T_229; // @[Shift.scala 90:48]
  wire [4:0] _GEN_7; // @[Shift.scala 90:39]
  wire [4:0] _T_231; // @[Shift.scala 90:39]
  wire  _T_233; // @[Shift.scala 12:21]
  wire [5:0] _T_234; // @[Cat.scala 29:58]
  wire [5:0] _T_235; // @[Shift.scala 91:22]
  wire [5:0] _T_238; // @[Bitwise.scala 71:12]
  wire [5:0] _T_239; // @[Shift.scala 39:10]
  wire  _T_240; // @[convert.scala 55:31]
  wire  _T_241; // @[convert.scala 56:31]
  wire  _T_242; // @[convert.scala 57:31]
  wire  _T_243; // @[convert.scala 58:31]
  wire [2:0] _T_244; // @[convert.scala 59:69]
  wire  _T_245; // @[convert.scala 59:81]
  wire  _T_246; // @[convert.scala 59:50]
  wire  _T_248; // @[convert.scala 60:81]
  wire  _T_249; // @[convert.scala 61:44]
  wire  _T_250; // @[convert.scala 61:52]
  wire  _T_251; // @[convert.scala 61:36]
  wire  _T_252; // @[convert.scala 62:63]
  wire  _T_253; // @[convert.scala 62:103]
  wire  _T_254; // @[convert.scala 62:60]
  wire [2:0] _GEN_8; // @[convert.scala 63:56]
  wire [2:0] _T_257; // @[convert.scala 63:56]
  wire [3:0] _T_258; // @[Cat.scala 29:58]
  reg  _T_262; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [3:0] _T_266; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  assign _T = io_quireIn[14:0]; // @[QuireToPosit.scala 47:43]
  assign _T_1 = _T != 15'h0; // @[QuireToPosit.scala 47:47]
  assign tailIsZero = ~ _T_1; // @[QuireToPosit.scala 47:27]
  assign _T_2 = io_quireIn[15:15]; // @[QuireToPosit.scala 49:45]
  assign outRawFloat_isNaR = _T_2 & tailIsZero; // @[QuireToPosit.scala 49:49]
  assign _T_5 = ~ _T_2; // @[QuireToPosit.scala 50:31]
  assign outRawFloat_isZero = _T_5 & tailIsZero; // @[QuireToPosit.scala 50:51]
  assign _T_8 = io_quireIn[15:1]; // @[QuireToPosit.scala 58:41]
  assign _T_9 = io_quireIn[14:0]; // @[QuireToPosit.scala 58:68]
  assign quireXOR = _T_8 ^ _T_9; // @[QuireToPosit.scala 58:56]
  assign _T_10 = quireXOR[14:7]; // @[LZD.scala 43:32]
  assign _T_11 = _T_10[7:4]; // @[LZD.scala 43:32]
  assign _T_12 = _T_11[3:2]; // @[LZD.scala 43:32]
  assign _T_13 = _T_12 != 2'h0; // @[LZD.scala 39:14]
  assign _T_14 = _T_12[1]; // @[LZD.scala 39:21]
  assign _T_15 = _T_12[0]; // @[LZD.scala 39:30]
  assign _T_16 = ~ _T_15; // @[LZD.scala 39:27]
  assign _T_17 = _T_14 | _T_16; // @[LZD.scala 39:25]
  assign _T_18 = {_T_13,_T_17}; // @[Cat.scala 29:58]
  assign _T_19 = _T_11[1:0]; // @[LZD.scala 44:32]
  assign _T_20 = _T_19 != 2'h0; // @[LZD.scala 39:14]
  assign _T_21 = _T_19[1]; // @[LZD.scala 39:21]
  assign _T_22 = _T_19[0]; // @[LZD.scala 39:30]
  assign _T_23 = ~ _T_22; // @[LZD.scala 39:27]
  assign _T_24 = _T_21 | _T_23; // @[LZD.scala 39:25]
  assign _T_25 = {_T_20,_T_24}; // @[Cat.scala 29:58]
  assign _T_26 = _T_18[1]; // @[Shift.scala 12:21]
  assign _T_27 = _T_25[1]; // @[Shift.scala 12:21]
  assign _T_28 = _T_26 | _T_27; // @[LZD.scala 49:16]
  assign _T_29 = ~ _T_27; // @[LZD.scala 49:27]
  assign _T_30 = _T_26 | _T_29; // @[LZD.scala 49:25]
  assign _T_31 = _T_18[0:0]; // @[LZD.scala 49:47]
  assign _T_32 = _T_25[0:0]; // @[LZD.scala 49:59]
  assign _T_33 = _T_26 ? _T_31 : _T_32; // @[LZD.scala 49:35]
  assign _T_35 = {_T_28,_T_30,_T_33}; // @[Cat.scala 29:58]
  assign _T_36 = _T_10[3:0]; // @[LZD.scala 44:32]
  assign _T_37 = _T_36[3:2]; // @[LZD.scala 43:32]
  assign _T_38 = _T_37 != 2'h0; // @[LZD.scala 39:14]
  assign _T_39 = _T_37[1]; // @[LZD.scala 39:21]
  assign _T_40 = _T_37[0]; // @[LZD.scala 39:30]
  assign _T_41 = ~ _T_40; // @[LZD.scala 39:27]
  assign _T_42 = _T_39 | _T_41; // @[LZD.scala 39:25]
  assign _T_43 = {_T_38,_T_42}; // @[Cat.scala 29:58]
  assign _T_44 = _T_36[1:0]; // @[LZD.scala 44:32]
  assign _T_45 = _T_44 != 2'h0; // @[LZD.scala 39:14]
  assign _T_46 = _T_44[1]; // @[LZD.scala 39:21]
  assign _T_47 = _T_44[0]; // @[LZD.scala 39:30]
  assign _T_48 = ~ _T_47; // @[LZD.scala 39:27]
  assign _T_49 = _T_46 | _T_48; // @[LZD.scala 39:25]
  assign _T_50 = {_T_45,_T_49}; // @[Cat.scala 29:58]
  assign _T_51 = _T_43[1]; // @[Shift.scala 12:21]
  assign _T_52 = _T_50[1]; // @[Shift.scala 12:21]
  assign _T_53 = _T_51 | _T_52; // @[LZD.scala 49:16]
  assign _T_54 = ~ _T_52; // @[LZD.scala 49:27]
  assign _T_55 = _T_51 | _T_54; // @[LZD.scala 49:25]
  assign _T_56 = _T_43[0:0]; // @[LZD.scala 49:47]
  assign _T_57 = _T_50[0:0]; // @[LZD.scala 49:59]
  assign _T_58 = _T_51 ? _T_56 : _T_57; // @[LZD.scala 49:35]
  assign _T_60 = {_T_53,_T_55,_T_58}; // @[Cat.scala 29:58]
  assign _T_61 = _T_35[2]; // @[Shift.scala 12:21]
  assign _T_62 = _T_60[2]; // @[Shift.scala 12:21]
  assign _T_63 = _T_61 | _T_62; // @[LZD.scala 49:16]
  assign _T_64 = ~ _T_62; // @[LZD.scala 49:27]
  assign _T_65 = _T_61 | _T_64; // @[LZD.scala 49:25]
  assign _T_66 = _T_35[1:0]; // @[LZD.scala 49:47]
  assign _T_67 = _T_60[1:0]; // @[LZD.scala 49:59]
  assign _T_68 = _T_61 ? _T_66 : _T_67; // @[LZD.scala 49:35]
  assign _T_70 = {_T_63,_T_65,_T_68}; // @[Cat.scala 29:58]
  assign _T_71 = quireXOR[6:0]; // @[LZD.scala 44:32]
  assign _T_72 = _T_71[6:3]; // @[LZD.scala 43:32]
  assign _T_73 = _T_72[3:2]; // @[LZD.scala 43:32]
  assign _T_74 = _T_73 != 2'h0; // @[LZD.scala 39:14]
  assign _T_75 = _T_73[1]; // @[LZD.scala 39:21]
  assign _T_76 = _T_73[0]; // @[LZD.scala 39:30]
  assign _T_77 = ~ _T_76; // @[LZD.scala 39:27]
  assign _T_78 = _T_75 | _T_77; // @[LZD.scala 39:25]
  assign _T_79 = {_T_74,_T_78}; // @[Cat.scala 29:58]
  assign _T_80 = _T_72[1:0]; // @[LZD.scala 44:32]
  assign _T_81 = _T_80 != 2'h0; // @[LZD.scala 39:14]
  assign _T_82 = _T_80[1]; // @[LZD.scala 39:21]
  assign _T_83 = _T_80[0]; // @[LZD.scala 39:30]
  assign _T_84 = ~ _T_83; // @[LZD.scala 39:27]
  assign _T_85 = _T_82 | _T_84; // @[LZD.scala 39:25]
  assign _T_86 = {_T_81,_T_85}; // @[Cat.scala 29:58]
  assign _T_87 = _T_79[1]; // @[Shift.scala 12:21]
  assign _T_88 = _T_86[1]; // @[Shift.scala 12:21]
  assign _T_89 = _T_87 | _T_88; // @[LZD.scala 49:16]
  assign _T_90 = ~ _T_88; // @[LZD.scala 49:27]
  assign _T_91 = _T_87 | _T_90; // @[LZD.scala 49:25]
  assign _T_92 = _T_79[0:0]; // @[LZD.scala 49:47]
  assign _T_93 = _T_86[0:0]; // @[LZD.scala 49:59]
  assign _T_94 = _T_87 ? _T_92 : _T_93; // @[LZD.scala 49:35]
  assign _T_96 = {_T_89,_T_91,_T_94}; // @[Cat.scala 29:58]
  assign _T_97 = _T_71[2:0]; // @[LZD.scala 44:32]
  assign _T_98 = _T_97[2:1]; // @[LZD.scala 43:32]
  assign _T_99 = _T_98 != 2'h0; // @[LZD.scala 39:14]
  assign _T_100 = _T_98[1]; // @[LZD.scala 39:21]
  assign _T_101 = _T_98[0]; // @[LZD.scala 39:30]
  assign _T_102 = ~ _T_101; // @[LZD.scala 39:27]
  assign _T_103 = _T_100 | _T_102; // @[LZD.scala 39:25]
  assign _T_104 = {_T_99,_T_103}; // @[Cat.scala 29:58]
  assign _T_105 = _T_97[0:0]; // @[LZD.scala 44:32]
  assign _T_107 = _T_104[1]; // @[Shift.scala 12:21]
  assign _T_109 = _T_104[0:0]; // @[LZD.scala 55:32]
  assign _T_110 = _T_107 ? _T_109 : _T_105; // @[LZD.scala 55:20]
  assign _T_111 = {_T_107,_T_110}; // @[Cat.scala 29:58]
  assign _T_112 = _T_96[2]; // @[Shift.scala 12:21]
  assign _T_114 = _T_96[1:0]; // @[LZD.scala 55:32]
  assign _T_115 = _T_112 ? _T_114 : _T_111; // @[LZD.scala 55:20]
  assign _T_116 = {_T_112,_T_115}; // @[Cat.scala 29:58]
  assign _T_117 = _T_70[3]; // @[Shift.scala 12:21]
  assign _T_119 = _T_70[2:0]; // @[LZD.scala 55:32]
  assign _T_120 = _T_117 ? _T_119 : _T_116; // @[LZD.scala 55:20]
  assign scaleBias = {1'h1,_T_117,_T_120}; // @[Cat.scala 29:58]
  assign _T_121 = $signed(scaleBias); // @[QuireToPosit.scala 61:53]
  assign _GEN_2 = {{1{_T_121[4]}},_T_121}; // @[QuireToPosit.scala 61:41]
  assign _T_123 = $signed(6'shb) + $signed(_GEN_2); // @[QuireToPosit.scala 61:41]
  assign realScale = $signed(_T_123); // @[QuireToPosit.scala 61:41]
  assign underflow = $signed(realScale) < $signed(-6'sh3); // @[QuireToPosit.scala 62:41]
  assign overflow = $signed(realScale) > $signed(6'sh2); // @[QuireToPosit.scala 63:35]
  assign _T_124 = underflow ? $signed(-6'sh3) : $signed(realScale); // @[Mux.scala 87:16]
  assign _T_125 = overflow ? $signed(6'sh2) : $signed(_T_124); // @[Mux.scala 87:16]
  assign _T_126 = realScale[5:5]; // @[Abs.scala 10:21]
  assign _T_128 = _T_126 ? 6'h3f : 6'h0; // @[Bitwise.scala 71:12]
  assign _T_129 = $unsigned(realScale); // @[Abs.scala 10:31]
  assign _T_130 = _T_128 ^ _T_129; // @[Abs.scala 10:26]
  assign _GEN_3 = {{5'd0}, _T_126}; // @[Abs.scala 10:39]
  assign absRealScale = _T_130 + _GEN_3; // @[Abs.scala 10:39]
  assign _T_133 = absRealScale < 6'h10; // @[Shift.scala 16:24]
  assign _T_134 = absRealScale[3:0]; // @[Shift.scala 17:37]
  assign _T_135 = _T_134[3]; // @[Shift.scala 12:21]
  assign _T_136 = io_quireIn[7:0]; // @[Shift.scala 64:52]
  assign _T_138 = {_T_136,8'h0}; // @[Cat.scala 29:58]
  assign _T_139 = _T_135 ? _T_138 : io_quireIn; // @[Shift.scala 64:27]
  assign _T_140 = _T_134[2:0]; // @[Shift.scala 66:70]
  assign _T_141 = _T_140[2]; // @[Shift.scala 12:21]
  assign _T_142 = _T_139[11:0]; // @[Shift.scala 64:52]
  assign _T_144 = {_T_142,4'h0}; // @[Cat.scala 29:58]
  assign _T_145 = _T_141 ? _T_144 : _T_139; // @[Shift.scala 64:27]
  assign _T_146 = _T_140[1:0]; // @[Shift.scala 66:70]
  assign _T_147 = _T_146[1]; // @[Shift.scala 12:21]
  assign _T_148 = _T_145[13:0]; // @[Shift.scala 64:52]
  assign _T_150 = {_T_148,2'h0}; // @[Cat.scala 29:58]
  assign _T_151 = _T_147 ? _T_150 : _T_145; // @[Shift.scala 64:27]
  assign _T_152 = _T_146[0:0]; // @[Shift.scala 66:70]
  assign _T_154 = _T_151[14:0]; // @[Shift.scala 64:52]
  assign _T_155 = {_T_154,1'h0}; // @[Cat.scala 29:58]
  assign _T_156 = _T_152 ? _T_155 : _T_151; // @[Shift.scala 64:27]
  assign quireLeftShift = _T_133 ? _T_156 : 16'h0; // @[Shift.scala 16:10]
  assign _T_161 = io_quireIn[15:8]; // @[Shift.scala 77:66]
  assign _T_162 = {8'h0,_T_161}; // @[Cat.scala 29:58]
  assign _T_163 = _T_135 ? _T_162 : io_quireIn; // @[Shift.scala 77:22]
  assign _T_167 = _T_163[15:4]; // @[Shift.scala 77:66]
  assign _T_168 = {4'h0,_T_167}; // @[Cat.scala 29:58]
  assign _T_169 = _T_141 ? _T_168 : _T_163; // @[Shift.scala 77:22]
  assign _T_173 = _T_169[15:2]; // @[Shift.scala 77:66]
  assign _T_174 = {2'h0,_T_173}; // @[Cat.scala 29:58]
  assign _T_175 = _T_147 ? _T_174 : _T_169; // @[Shift.scala 77:22]
  assign _T_178 = _T_175[15:1]; // @[Shift.scala 77:66]
  assign _T_179 = {1'h0,_T_178}; // @[Cat.scala 29:58]
  assign _T_180 = _T_152 ? _T_179 : _T_175; // @[Shift.scala 77:22]
  assign quireRightShift = _T_133 ? _T_180 : 16'h0; // @[Shift.scala 27:10]
  assign _T_182 = quireLeftShift[3:1]; // @[QuireToPosit.scala 89:49]
  assign _T_183 = quireLeftShift[0]; // @[QuireToPosit.scala 90:127]
  assign realFGRSTmp1 = {_T_182,_T_183}; // @[Cat.scala 29:58]
  assign _T_185 = quireRightShift[3:1]; // @[QuireToPosit.scala 91:50]
  assign _T_186 = quireRightShift[0]; // @[QuireToPosit.scala 92:128]
  assign realFGRSTmp2 = {_T_185,_T_186}; // @[Cat.scala 29:58]
  assign realFGRS = _T_126 ? realFGRSTmp1 : realFGRSTmp2; // @[QuireToPosit.scala 93:34]
  assign outRawFloat_fraction = realFGRS[3:3]; // @[QuireToPosit.scala 95:46]
  assign outRawFloat_grs = realFGRS[2:0]; // @[QuireToPosit.scala 96:46]
  assign _GEN_4 = _T_125[2:0]; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  assign outRawFloat_scale = $signed(_GEN_4); // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  assign _T_193 = outRawFloat_scale[2:2]; // @[convert.scala 49:36]
  assign _T_195 = ~ outRawFloat_scale; // @[convert.scala 50:36]
  assign _T_196 = $signed(_T_195); // @[convert.scala 50:36]
  assign _T_197 = _T_193 ? $signed(_T_196) : $signed(outRawFloat_scale); // @[convert.scala 50:28]
  assign _T_198 = _T_193 ^ _T_2; // @[convert.scala 51:31]
  assign _T_199 = ~ _T_198; // @[convert.scala 53:34]
  assign _T_202 = {_T_199,_T_198,outRawFloat_fraction,outRawFloat_grs}; // @[Cat.scala 29:58]
  assign _T_203 = $unsigned(_T_197); // @[Shift.scala 39:17]
  assign _T_204 = _T_203 < 3'h6; // @[Shift.scala 39:24]
  assign _T_206 = _T_202[5:4]; // @[Shift.scala 90:30]
  assign _T_207 = _T_202[3:0]; // @[Shift.scala 90:48]
  assign _T_208 = _T_207 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{1'd0}, _T_208}; // @[Shift.scala 90:39]
  assign _T_209 = _T_206 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_210 = _T_203[2]; // @[Shift.scala 12:21]
  assign _T_211 = _T_202[5]; // @[Shift.scala 12:21]
  assign _T_213 = _T_211 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_214 = {_T_213,_T_209}; // @[Cat.scala 29:58]
  assign _T_215 = _T_210 ? _T_214 : _T_202; // @[Shift.scala 91:22]
  assign _T_216 = _T_203[1:0]; // @[Shift.scala 92:77]
  assign _T_217 = _T_215[5:2]; // @[Shift.scala 90:30]
  assign _T_218 = _T_215[1:0]; // @[Shift.scala 90:48]
  assign _T_219 = _T_218 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{3'd0}, _T_219}; // @[Shift.scala 90:39]
  assign _T_220 = _T_217 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_221 = _T_216[1]; // @[Shift.scala 12:21]
  assign _T_222 = _T_215[5]; // @[Shift.scala 12:21]
  assign _T_224 = _T_222 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_225 = {_T_224,_T_220}; // @[Cat.scala 29:58]
  assign _T_226 = _T_221 ? _T_225 : _T_215; // @[Shift.scala 91:22]
  assign _T_227 = _T_216[0:0]; // @[Shift.scala 92:77]
  assign _T_228 = _T_226[5:1]; // @[Shift.scala 90:30]
  assign _T_229 = _T_226[0:0]; // @[Shift.scala 90:48]
  assign _GEN_7 = {{4'd0}, _T_229}; // @[Shift.scala 90:39]
  assign _T_231 = _T_228 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_233 = _T_226[5]; // @[Shift.scala 12:21]
  assign _T_234 = {_T_233,_T_231}; // @[Cat.scala 29:58]
  assign _T_235 = _T_227 ? _T_234 : _T_226; // @[Shift.scala 91:22]
  assign _T_238 = _T_211 ? 6'h3f : 6'h0; // @[Bitwise.scala 71:12]
  assign _T_239 = _T_204 ? _T_235 : _T_238; // @[Shift.scala 39:10]
  assign _T_240 = _T_239[3]; // @[convert.scala 55:31]
  assign _T_241 = _T_239[2]; // @[convert.scala 56:31]
  assign _T_242 = _T_239[1]; // @[convert.scala 57:31]
  assign _T_243 = _T_239[0]; // @[convert.scala 58:31]
  assign _T_244 = _T_239[5:3]; // @[convert.scala 59:69]
  assign _T_245 = _T_244 != 3'h0; // @[convert.scala 59:81]
  assign _T_246 = ~ _T_245; // @[convert.scala 59:50]
  assign _T_248 = _T_244 == 3'h7; // @[convert.scala 60:81]
  assign _T_249 = _T_240 | _T_242; // @[convert.scala 61:44]
  assign _T_250 = _T_249 | _T_243; // @[convert.scala 61:52]
  assign _T_251 = _T_241 & _T_250; // @[convert.scala 61:36]
  assign _T_252 = ~ _T_248; // @[convert.scala 62:63]
  assign _T_253 = _T_252 & _T_251; // @[convert.scala 62:103]
  assign _T_254 = _T_246 | _T_253; // @[convert.scala 62:60]
  assign _GEN_8 = {{2'd0}, _T_254}; // @[convert.scala 63:56]
  assign _T_257 = _T_244 + _GEN_8; // @[convert.scala 63:56]
  assign _T_258 = {_T_2,_T_257}; // @[Cat.scala 29:58]
  assign io_positOut = _T_266; // @[QuireToPosit.scala 101:15]
  assign io_outValid = _T_262; // @[QuireToPosit.scala 100:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_262 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_266 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_262 <= 1'h0;
    end else begin
      _T_262 <= io_inValid;
    end
    if (io_inValid) begin
      if (outRawFloat_isNaR) begin
        _T_266 <= 4'h8;
      end else begin
        if (outRawFloat_isZero) begin
          _T_266 <= 4'h0;
        end else begin
          _T_266 <= _T_258;
        end
      end
    end
  end
endmodule
