module PositFMA6_0(
  input        clock,
  input        reset,
  input        io_inValid,
  input  [1:0] io_fmaOp,
  input  [5:0] io_A,
  input  [5:0] io_B,
  input  [5:0] io_C,
  output [5:0] io_F,
  output       io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [5:0] _T_2; // @[Bitwise.scala 71:12]
  wire [5:0] _T_3; // @[PositFMA.scala 47:41]
  wire [5:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [5:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [5:0] _T_8; // @[Bitwise.scala 71:12]
  wire [5:0] _T_9; // @[PositFMA.scala 48:41]
  wire [5:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [5:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [3:0] _T_16; // @[convert.scala 19:24]
  wire [3:0] _T_17; // @[convert.scala 19:43]
  wire [3:0] _T_18; // @[convert.scala 19:39]
  wire [1:0] _T_19; // @[LZD.scala 43:32]
  wire  _T_20; // @[LZD.scala 39:14]
  wire  _T_21; // @[LZD.scala 39:21]
  wire  _T_22; // @[LZD.scala 39:30]
  wire  _T_23; // @[LZD.scala 39:27]
  wire  _T_24; // @[LZD.scala 39:25]
  wire [1:0] _T_25; // @[Cat.scala 29:58]
  wire [1:0] _T_26; // @[LZD.scala 44:32]
  wire  _T_27; // @[LZD.scala 39:14]
  wire  _T_28; // @[LZD.scala 39:21]
  wire  _T_29; // @[LZD.scala 39:30]
  wire  _T_30; // @[LZD.scala 39:27]
  wire  _T_31; // @[LZD.scala 39:25]
  wire [1:0] _T_32; // @[Cat.scala 29:58]
  wire  _T_33; // @[Shift.scala 12:21]
  wire  _T_34; // @[Shift.scala 12:21]
  wire  _T_35; // @[LZD.scala 49:16]
  wire  _T_36; // @[LZD.scala 49:27]
  wire  _T_37; // @[LZD.scala 49:25]
  wire  _T_38; // @[LZD.scala 49:47]
  wire  _T_39; // @[LZD.scala 49:59]
  wire  _T_40; // @[LZD.scala 49:35]
  wire [2:0] _T_42; // @[Cat.scala 29:58]
  wire [2:0] _T_43; // @[convert.scala 21:22]
  wire [2:0] _T_44; // @[convert.scala 22:36]
  wire  _T_45; // @[Shift.scala 16:24]
  wire [1:0] _T_46; // @[Shift.scala 17:37]
  wire  _T_47; // @[Shift.scala 12:21]
  wire  _T_48; // @[Shift.scala 64:52]
  wire [2:0] _T_50; // @[Cat.scala 29:58]
  wire [2:0] _T_51; // @[Shift.scala 64:27]
  wire  _T_52; // @[Shift.scala 66:70]
  wire [1:0] _T_54; // @[Shift.scala 64:52]
  wire [2:0] _T_55; // @[Cat.scala 29:58]
  wire [2:0] _T_56; // @[Shift.scala 64:27]
  wire [2:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_60; // @[convert.scala 25:26]
  wire [2:0] _T_62; // @[convert.scala 25:42]
  wire [3:0] _T_63; // @[Cat.scala 29:58]
  wire [4:0] _T_65; // @[convert.scala 29:56]
  wire  _T_66; // @[convert.scala 29:60]
  wire  _T_67; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_70; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [3:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_79; // @[convert.scala 18:24]
  wire  _T_80; // @[convert.scala 18:40]
  wire  _T_81; // @[convert.scala 18:36]
  wire [3:0] _T_82; // @[convert.scala 19:24]
  wire [3:0] _T_83; // @[convert.scala 19:43]
  wire [3:0] _T_84; // @[convert.scala 19:39]
  wire [1:0] _T_85; // @[LZD.scala 43:32]
  wire  _T_86; // @[LZD.scala 39:14]
  wire  _T_87; // @[LZD.scala 39:21]
  wire  _T_88; // @[LZD.scala 39:30]
  wire  _T_89; // @[LZD.scala 39:27]
  wire  _T_90; // @[LZD.scala 39:25]
  wire [1:0] _T_91; // @[Cat.scala 29:58]
  wire [1:0] _T_92; // @[LZD.scala 44:32]
  wire  _T_93; // @[LZD.scala 39:14]
  wire  _T_94; // @[LZD.scala 39:21]
  wire  _T_95; // @[LZD.scala 39:30]
  wire  _T_96; // @[LZD.scala 39:27]
  wire  _T_97; // @[LZD.scala 39:25]
  wire [1:0] _T_98; // @[Cat.scala 29:58]
  wire  _T_99; // @[Shift.scala 12:21]
  wire  _T_100; // @[Shift.scala 12:21]
  wire  _T_101; // @[LZD.scala 49:16]
  wire  _T_102; // @[LZD.scala 49:27]
  wire  _T_103; // @[LZD.scala 49:25]
  wire  _T_104; // @[LZD.scala 49:47]
  wire  _T_105; // @[LZD.scala 49:59]
  wire  _T_106; // @[LZD.scala 49:35]
  wire [2:0] _T_108; // @[Cat.scala 29:58]
  wire [2:0] _T_109; // @[convert.scala 21:22]
  wire [2:0] _T_110; // @[convert.scala 22:36]
  wire  _T_111; // @[Shift.scala 16:24]
  wire [1:0] _T_112; // @[Shift.scala 17:37]
  wire  _T_113; // @[Shift.scala 12:21]
  wire  _T_114; // @[Shift.scala 64:52]
  wire [2:0] _T_116; // @[Cat.scala 29:58]
  wire [2:0] _T_117; // @[Shift.scala 64:27]
  wire  _T_118; // @[Shift.scala 66:70]
  wire [1:0] _T_120; // @[Shift.scala 64:52]
  wire [2:0] _T_121; // @[Cat.scala 29:58]
  wire [2:0] _T_122; // @[Shift.scala 64:27]
  wire [2:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_126; // @[convert.scala 25:26]
  wire [2:0] _T_128; // @[convert.scala 25:42]
  wire [3:0] _T_129; // @[Cat.scala 29:58]
  wire [4:0] _T_131; // @[convert.scala 29:56]
  wire  _T_132; // @[convert.scala 29:60]
  wire  _T_133; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_136; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [3:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_145; // @[convert.scala 18:24]
  wire  _T_146; // @[convert.scala 18:40]
  wire  _T_147; // @[convert.scala 18:36]
  wire [3:0] _T_148; // @[convert.scala 19:24]
  wire [3:0] _T_149; // @[convert.scala 19:43]
  wire [3:0] _T_150; // @[convert.scala 19:39]
  wire [1:0] _T_151; // @[LZD.scala 43:32]
  wire  _T_152; // @[LZD.scala 39:14]
  wire  _T_153; // @[LZD.scala 39:21]
  wire  _T_154; // @[LZD.scala 39:30]
  wire  _T_155; // @[LZD.scala 39:27]
  wire  _T_156; // @[LZD.scala 39:25]
  wire [1:0] _T_157; // @[Cat.scala 29:58]
  wire [1:0] _T_158; // @[LZD.scala 44:32]
  wire  _T_159; // @[LZD.scala 39:14]
  wire  _T_160; // @[LZD.scala 39:21]
  wire  _T_161; // @[LZD.scala 39:30]
  wire  _T_162; // @[LZD.scala 39:27]
  wire  _T_163; // @[LZD.scala 39:25]
  wire [1:0] _T_164; // @[Cat.scala 29:58]
  wire  _T_165; // @[Shift.scala 12:21]
  wire  _T_166; // @[Shift.scala 12:21]
  wire  _T_167; // @[LZD.scala 49:16]
  wire  _T_168; // @[LZD.scala 49:27]
  wire  _T_169; // @[LZD.scala 49:25]
  wire  _T_170; // @[LZD.scala 49:47]
  wire  _T_171; // @[LZD.scala 49:59]
  wire  _T_172; // @[LZD.scala 49:35]
  wire [2:0] _T_174; // @[Cat.scala 29:58]
  wire [2:0] _T_175; // @[convert.scala 21:22]
  wire [2:0] _T_176; // @[convert.scala 22:36]
  wire  _T_177; // @[Shift.scala 16:24]
  wire [1:0] _T_178; // @[Shift.scala 17:37]
  wire  _T_179; // @[Shift.scala 12:21]
  wire  _T_180; // @[Shift.scala 64:52]
  wire [2:0] _T_182; // @[Cat.scala 29:58]
  wire [2:0] _T_183; // @[Shift.scala 64:27]
  wire  _T_184; // @[Shift.scala 66:70]
  wire [1:0] _T_186; // @[Shift.scala 64:52]
  wire [2:0] _T_187; // @[Cat.scala 29:58]
  wire  _T_192; // @[convert.scala 25:26]
  wire [2:0] _T_194; // @[convert.scala 25:42]
  wire [3:0] _T_195; // @[Cat.scala 29:58]
  wire [4:0] _T_197; // @[convert.scala 29:56]
  wire  _T_198; // @[convert.scala 29:60]
  wire  _T_199; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_202; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [3:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_210; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_211; // @[PositFMA.scala 59:34]
  wire  _T_212; // @[PositFMA.scala 59:47]
  wire  _T_213; // @[PositFMA.scala 59:45]
  wire [4:0] _T_215; // @[Cat.scala 29:58]
  wire [4:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_216; // @[PositFMA.scala 60:34]
  wire  _T_217; // @[PositFMA.scala 60:47]
  wire  _T_218; // @[PositFMA.scala 60:45]
  wire [4:0] _T_220; // @[Cat.scala 29:58]
  wire [4:0] sigB; // @[PositFMA.scala 60:76]
  wire [9:0] _T_221; // @[PositFMA.scala 62:25]
  wire [9:0] sigP; // @[PositFMA.scala 62:33]
  wire [1:0] head2; // @[PositFMA.scala 63:28]
  wire  _T_222; // @[PositFMA.scala 64:31]
  wire  _T_223; // @[PositFMA.scala 64:25]
  wire  _T_224; // @[PositFMA.scala 64:42]
  wire  addTwo; // @[PositFMA.scala 64:35]
  wire  _T_225; // @[PositFMA.scala 66:23]
  wire  _T_226; // @[PositFMA.scala 66:49]
  wire  addOne; // @[PositFMA.scala 66:43]
  wire [1:0] _T_227; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 67:39]
  wire  mulSign; // @[PositFMA.scala 68:28]
  wire [4:0] _T_228; // @[PositFMA.scala 70:30]
  wire [4:0] _GEN_12; // @[PositFMA.scala 70:44]
  wire [4:0] _T_230; // @[PositFMA.scala 70:44]
  wire [4:0] mulScale; // @[PositFMA.scala 70:44]
  wire [7:0] _T_231; // @[PositFMA.scala 73:29]
  wire [6:0] _T_232; // @[PositFMA.scala 74:29]
  wire [7:0] _T_233; // @[PositFMA.scala 74:48]
  wire [7:0] mulSigTmp; // @[PositFMA.scala 71:22]
  wire  _T_235; // @[PositFMA.scala 78:39]
  wire  _T_236; // @[PositFMA.scala 78:43]
  wire [6:0] _T_237; // @[PositFMA.scala 79:39]
  wire [8:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [8:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [2:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [4:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [3:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_263; // @[PositFMA.scala 108:29]
  wire  _T_264; // @[PositFMA.scala 108:47]
  wire  _T_265; // @[PositFMA.scala 108:45]
  wire [8:0] extAddSig; // @[Cat.scala 29:58]
  wire [4:0] _GEN_13; // @[PositFMA.scala 112:39]
  wire  mulGreater; // @[PositFMA.scala 112:39]
  wire [4:0] greaterScale; // @[PositFMA.scala 113:26]
  wire [4:0] smallerScale; // @[PositFMA.scala 114:26]
  wire [4:0] _T_269; // @[PositFMA.scala 115:36]
  wire [4:0] scaleDiff; // @[PositFMA.scala 115:36]
  wire [8:0] greaterSig; // @[PositFMA.scala 116:26]
  wire [8:0] smallerSigTmp; // @[PositFMA.scala 117:26]
  wire [4:0] _T_270; // @[PositFMA.scala 118:69]
  wire  _T_271; // @[Shift.scala 39:24]
  wire [3:0] _T_272; // @[Shift.scala 40:44]
  wire  _T_273; // @[Shift.scala 90:30]
  wire [7:0] _T_274; // @[Shift.scala 90:48]
  wire  _T_275; // @[Shift.scala 90:57]
  wire  _T_276; // @[Shift.scala 90:39]
  wire  _T_277; // @[Shift.scala 12:21]
  wire  _T_278; // @[Shift.scala 12:21]
  wire [7:0] _T_280; // @[Bitwise.scala 71:12]
  wire [8:0] _T_281; // @[Cat.scala 29:58]
  wire [8:0] _T_282; // @[Shift.scala 91:22]
  wire [2:0] _T_283; // @[Shift.scala 92:77]
  wire [4:0] _T_284; // @[Shift.scala 90:30]
  wire [3:0] _T_285; // @[Shift.scala 90:48]
  wire  _T_286; // @[Shift.scala 90:57]
  wire [4:0] _GEN_14; // @[Shift.scala 90:39]
  wire [4:0] _T_287; // @[Shift.scala 90:39]
  wire  _T_288; // @[Shift.scala 12:21]
  wire  _T_289; // @[Shift.scala 12:21]
  wire [3:0] _T_291; // @[Bitwise.scala 71:12]
  wire [8:0] _T_292; // @[Cat.scala 29:58]
  wire [8:0] _T_293; // @[Shift.scala 91:22]
  wire [1:0] _T_294; // @[Shift.scala 92:77]
  wire [6:0] _T_295; // @[Shift.scala 90:30]
  wire [1:0] _T_296; // @[Shift.scala 90:48]
  wire  _T_297; // @[Shift.scala 90:57]
  wire [6:0] _GEN_15; // @[Shift.scala 90:39]
  wire [6:0] _T_298; // @[Shift.scala 90:39]
  wire  _T_299; // @[Shift.scala 12:21]
  wire  _T_300; // @[Shift.scala 12:21]
  wire [1:0] _T_302; // @[Bitwise.scala 71:12]
  wire [8:0] _T_303; // @[Cat.scala 29:58]
  wire [8:0] _T_304; // @[Shift.scala 91:22]
  wire  _T_305; // @[Shift.scala 92:77]
  wire [7:0] _T_306; // @[Shift.scala 90:30]
  wire  _T_307; // @[Shift.scala 90:48]
  wire [7:0] _GEN_16; // @[Shift.scala 90:39]
  wire [7:0] _T_309; // @[Shift.scala 90:39]
  wire  _T_311; // @[Shift.scala 12:21]
  wire [8:0] _T_312; // @[Cat.scala 29:58]
  wire [8:0] _T_313; // @[Shift.scala 91:22]
  wire [8:0] _T_316; // @[Bitwise.scala 71:12]
  wire [8:0] smallerSig; // @[Shift.scala 39:10]
  wire [9:0] rawSumSig; // @[PositFMA.scala 119:34]
  wire  _T_317; // @[PositFMA.scala 120:42]
  wire  _T_318; // @[PositFMA.scala 120:46]
  wire  _T_319; // @[PositFMA.scala 120:79]
  wire  sumSign; // @[PositFMA.scala 120:63]
  wire [8:0] _T_321; // @[PositFMA.scala 121:50]
  wire [9:0] signSumSig; // @[Cat.scala 29:58]
  wire [8:0] _T_322; // @[PositFMA.scala 126:33]
  wire [8:0] _T_323; // @[PositFMA.scala 126:68]
  wire [8:0] sumXor; // @[PositFMA.scala 126:51]
  wire [7:0] _T_324; // @[LZD.scala 43:32]
  wire [3:0] _T_325; // @[LZD.scala 43:32]
  wire [1:0] _T_326; // @[LZD.scala 43:32]
  wire  _T_327; // @[LZD.scala 39:14]
  wire  _T_328; // @[LZD.scala 39:21]
  wire  _T_329; // @[LZD.scala 39:30]
  wire  _T_330; // @[LZD.scala 39:27]
  wire  _T_331; // @[LZD.scala 39:25]
  wire [1:0] _T_332; // @[Cat.scala 29:58]
  wire [1:0] _T_333; // @[LZD.scala 44:32]
  wire  _T_334; // @[LZD.scala 39:14]
  wire  _T_335; // @[LZD.scala 39:21]
  wire  _T_336; // @[LZD.scala 39:30]
  wire  _T_337; // @[LZD.scala 39:27]
  wire  _T_338; // @[LZD.scala 39:25]
  wire [1:0] _T_339; // @[Cat.scala 29:58]
  wire  _T_340; // @[Shift.scala 12:21]
  wire  _T_341; // @[Shift.scala 12:21]
  wire  _T_342; // @[LZD.scala 49:16]
  wire  _T_343; // @[LZD.scala 49:27]
  wire  _T_344; // @[LZD.scala 49:25]
  wire  _T_345; // @[LZD.scala 49:47]
  wire  _T_346; // @[LZD.scala 49:59]
  wire  _T_347; // @[LZD.scala 49:35]
  wire [2:0] _T_349; // @[Cat.scala 29:58]
  wire [3:0] _T_350; // @[LZD.scala 44:32]
  wire [1:0] _T_351; // @[LZD.scala 43:32]
  wire  _T_352; // @[LZD.scala 39:14]
  wire  _T_353; // @[LZD.scala 39:21]
  wire  _T_354; // @[LZD.scala 39:30]
  wire  _T_355; // @[LZD.scala 39:27]
  wire  _T_356; // @[LZD.scala 39:25]
  wire [1:0] _T_357; // @[Cat.scala 29:58]
  wire [1:0] _T_358; // @[LZD.scala 44:32]
  wire  _T_359; // @[LZD.scala 39:14]
  wire  _T_360; // @[LZD.scala 39:21]
  wire  _T_361; // @[LZD.scala 39:30]
  wire  _T_362; // @[LZD.scala 39:27]
  wire  _T_363; // @[LZD.scala 39:25]
  wire [1:0] _T_364; // @[Cat.scala 29:58]
  wire  _T_365; // @[Shift.scala 12:21]
  wire  _T_366; // @[Shift.scala 12:21]
  wire  _T_367; // @[LZD.scala 49:16]
  wire  _T_368; // @[LZD.scala 49:27]
  wire  _T_369; // @[LZD.scala 49:25]
  wire  _T_370; // @[LZD.scala 49:47]
  wire  _T_371; // @[LZD.scala 49:59]
  wire  _T_372; // @[LZD.scala 49:35]
  wire [2:0] _T_374; // @[Cat.scala 29:58]
  wire  _T_375; // @[Shift.scala 12:21]
  wire  _T_376; // @[Shift.scala 12:21]
  wire  _T_377; // @[LZD.scala 49:16]
  wire  _T_378; // @[LZD.scala 49:27]
  wire  _T_379; // @[LZD.scala 49:25]
  wire [1:0] _T_380; // @[LZD.scala 49:47]
  wire [1:0] _T_381; // @[LZD.scala 49:59]
  wire [1:0] _T_382; // @[LZD.scala 49:35]
  wire [3:0] _T_384; // @[Cat.scala 29:58]
  wire  _T_385; // @[LZD.scala 44:32]
  wire  _T_387; // @[Shift.scala 12:21]
  wire [2:0] _T_390; // @[Cat.scala 29:58]
  wire [2:0] _T_391; // @[LZD.scala 55:32]
  wire [2:0] _T_392; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [3:0] shiftValue; // @[PositFMA.scala 128:24]
  wire [7:0] _T_393; // @[PositFMA.scala 129:38]
  wire  _T_394; // @[Shift.scala 16:24]
  wire [2:0] _T_395; // @[Shift.scala 17:37]
  wire  _T_396; // @[Shift.scala 12:21]
  wire [3:0] _T_397; // @[Shift.scala 64:52]
  wire [7:0] _T_399; // @[Cat.scala 29:58]
  wire [7:0] _T_400; // @[Shift.scala 64:27]
  wire [1:0] _T_401; // @[Shift.scala 66:70]
  wire  _T_402; // @[Shift.scala 12:21]
  wire [5:0] _T_403; // @[Shift.scala 64:52]
  wire [7:0] _T_405; // @[Cat.scala 29:58]
  wire [7:0] _T_406; // @[Shift.scala 64:27]
  wire  _T_407; // @[Shift.scala 66:70]
  wire [6:0] _T_409; // @[Shift.scala 64:52]
  wire [7:0] _T_410; // @[Cat.scala 29:58]
  wire [7:0] _T_411; // @[Shift.scala 64:27]
  wire [7:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [4:0] _T_413; // @[PositFMA.scala 132:36]
  wire [4:0] _T_414; // @[PositFMA.scala 132:36]
  wire [4:0] _T_415; // @[Cat.scala 29:58]
  wire [4:0] _T_416; // @[PositFMA.scala 132:61]
  wire [4:0] _T_418; // @[PositFMA.scala 132:42]
  wire [4:0] sumScale; // @[PositFMA.scala 132:42]
  wire [2:0] sumFrac; // @[PositFMA.scala 133:41]
  wire [4:0] grsTmp; // @[PositFMA.scala 136:41]
  wire [1:0] _T_419; // @[PositFMA.scala 139:40]
  wire [2:0] _T_420; // @[PositFMA.scala 139:56]
  wire  _T_421; // @[PositFMA.scala 139:60]
  wire  underflow; // @[PositFMA.scala 146:32]
  wire  overflow; // @[PositFMA.scala 147:32]
  wire  _T_422; // @[PositFMA.scala 156:32]
  wire  decF_isZero; // @[PositFMA.scala 156:20]
  wire [4:0] _T_424; // @[Mux.scala 87:16]
  wire [4:0] _T_425; // @[Mux.scala 87:16]
  wire [3:0] _GEN_17; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  wire [3:0] decF_scale; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  wire  _T_427; // @[convert.scala 49:36]
  wire [3:0] _T_429; // @[convert.scala 50:36]
  wire [3:0] _T_430; // @[convert.scala 50:36]
  wire [3:0] _T_431; // @[convert.scala 50:28]
  wire  _T_432; // @[convert.scala 51:31]
  wire  _T_433; // @[convert.scala 53:34]
  wire [7:0] _T_436; // @[Cat.scala 29:58]
  wire [3:0] _T_437; // @[Shift.scala 39:17]
  wire  _T_438; // @[Shift.scala 39:24]
  wire [2:0] _T_439; // @[Shift.scala 40:44]
  wire [3:0] _T_440; // @[Shift.scala 90:30]
  wire [3:0] _T_441; // @[Shift.scala 90:48]
  wire  _T_442; // @[Shift.scala 90:57]
  wire [3:0] _GEN_18; // @[Shift.scala 90:39]
  wire [3:0] _T_443; // @[Shift.scala 90:39]
  wire  _T_444; // @[Shift.scala 12:21]
  wire  _T_445; // @[Shift.scala 12:21]
  wire [3:0] _T_447; // @[Bitwise.scala 71:12]
  wire [7:0] _T_448; // @[Cat.scala 29:58]
  wire [7:0] _T_449; // @[Shift.scala 91:22]
  wire [1:0] _T_450; // @[Shift.scala 92:77]
  wire [5:0] _T_451; // @[Shift.scala 90:30]
  wire [1:0] _T_452; // @[Shift.scala 90:48]
  wire  _T_453; // @[Shift.scala 90:57]
  wire [5:0] _GEN_19; // @[Shift.scala 90:39]
  wire [5:0] _T_454; // @[Shift.scala 90:39]
  wire  _T_455; // @[Shift.scala 12:21]
  wire  _T_456; // @[Shift.scala 12:21]
  wire [1:0] _T_458; // @[Bitwise.scala 71:12]
  wire [7:0] _T_459; // @[Cat.scala 29:58]
  wire [7:0] _T_460; // @[Shift.scala 91:22]
  wire  _T_461; // @[Shift.scala 92:77]
  wire [6:0] _T_462; // @[Shift.scala 90:30]
  wire  _T_463; // @[Shift.scala 90:48]
  wire [6:0] _GEN_20; // @[Shift.scala 90:39]
  wire [6:0] _T_465; // @[Shift.scala 90:39]
  wire  _T_467; // @[Shift.scala 12:21]
  wire [7:0] _T_468; // @[Cat.scala 29:58]
  wire [7:0] _T_469; // @[Shift.scala 91:22]
  wire [7:0] _T_472; // @[Bitwise.scala 71:12]
  wire [7:0] _T_473; // @[Shift.scala 39:10]
  wire  _T_474; // @[convert.scala 55:31]
  wire  _T_475; // @[convert.scala 56:31]
  wire  _T_476; // @[convert.scala 57:31]
  wire  _T_477; // @[convert.scala 58:31]
  wire [4:0] _T_478; // @[convert.scala 59:69]
  wire  _T_479; // @[convert.scala 59:81]
  wire  _T_480; // @[convert.scala 59:50]
  wire  _T_482; // @[convert.scala 60:81]
  wire  _T_483; // @[convert.scala 61:44]
  wire  _T_484; // @[convert.scala 61:52]
  wire  _T_485; // @[convert.scala 61:36]
  wire  _T_486; // @[convert.scala 62:63]
  wire  _T_487; // @[convert.scala 62:103]
  wire  _T_488; // @[convert.scala 62:60]
  wire [4:0] _GEN_21; // @[convert.scala 63:56]
  wire [4:0] _T_491; // @[convert.scala 63:56]
  wire [5:0] _T_492; // @[Cat.scala 29:58]
  reg  _T_496; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [5:0] _T_500; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 6'h3f : 6'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{5'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 6'h3f : 6'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{5'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[5]; // @[convert.scala 18:24]
  assign _T_14 = realA[4]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[4:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[3:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[3:2]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19 != 2'h0; // @[LZD.scala 39:14]
  assign _T_21 = _T_19[1]; // @[LZD.scala 39:21]
  assign _T_22 = _T_19[0]; // @[LZD.scala 39:30]
  assign _T_23 = ~ _T_22; // @[LZD.scala 39:27]
  assign _T_24 = _T_21 | _T_23; // @[LZD.scala 39:25]
  assign _T_25 = {_T_20,_T_24}; // @[Cat.scala 29:58]
  assign _T_26 = _T_18[1:0]; // @[LZD.scala 44:32]
  assign _T_27 = _T_26 != 2'h0; // @[LZD.scala 39:14]
  assign _T_28 = _T_26[1]; // @[LZD.scala 39:21]
  assign _T_29 = _T_26[0]; // @[LZD.scala 39:30]
  assign _T_30 = ~ _T_29; // @[LZD.scala 39:27]
  assign _T_31 = _T_28 | _T_30; // @[LZD.scala 39:25]
  assign _T_32 = {_T_27,_T_31}; // @[Cat.scala 29:58]
  assign _T_33 = _T_25[1]; // @[Shift.scala 12:21]
  assign _T_34 = _T_32[1]; // @[Shift.scala 12:21]
  assign _T_35 = _T_33 | _T_34; // @[LZD.scala 49:16]
  assign _T_36 = ~ _T_34; // @[LZD.scala 49:27]
  assign _T_37 = _T_33 | _T_36; // @[LZD.scala 49:25]
  assign _T_38 = _T_25[0:0]; // @[LZD.scala 49:47]
  assign _T_39 = _T_32[0:0]; // @[LZD.scala 49:59]
  assign _T_40 = _T_33 ? _T_38 : _T_39; // @[LZD.scala 49:35]
  assign _T_42 = {_T_35,_T_37,_T_40}; // @[Cat.scala 29:58]
  assign _T_43 = ~ _T_42; // @[convert.scala 21:22]
  assign _T_44 = realA[2:0]; // @[convert.scala 22:36]
  assign _T_45 = _T_43 < 3'h3; // @[Shift.scala 16:24]
  assign _T_46 = _T_43[1:0]; // @[Shift.scala 17:37]
  assign _T_47 = _T_46[1]; // @[Shift.scala 12:21]
  assign _T_48 = _T_44[0:0]; // @[Shift.scala 64:52]
  assign _T_50 = {_T_48,2'h0}; // @[Cat.scala 29:58]
  assign _T_51 = _T_47 ? _T_50 : _T_44; // @[Shift.scala 64:27]
  assign _T_52 = _T_46[0:0]; // @[Shift.scala 66:70]
  assign _T_54 = _T_51[1:0]; // @[Shift.scala 64:52]
  assign _T_55 = {_T_54,1'h0}; // @[Cat.scala 29:58]
  assign _T_56 = _T_52 ? _T_55 : _T_51; // @[Shift.scala 64:27]
  assign decA_fraction = _T_45 ? _T_56 : 3'h0; // @[Shift.scala 16:10]
  assign _T_60 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_62 = _T_15 ? _T_43 : _T_42; // @[convert.scala 25:42]
  assign _T_63 = {_T_60,_T_62}; // @[Cat.scala 29:58]
  assign _T_65 = realA[4:0]; // @[convert.scala 29:56]
  assign _T_66 = _T_65 != 5'h0; // @[convert.scala 29:60]
  assign _T_67 = ~ _T_66; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_67; // @[convert.scala 29:39]
  assign _T_70 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_70 & _T_67; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_63); // @[convert.scala 32:24]
  assign _T_79 = io_B[5]; // @[convert.scala 18:24]
  assign _T_80 = io_B[4]; // @[convert.scala 18:40]
  assign _T_81 = _T_79 ^ _T_80; // @[convert.scala 18:36]
  assign _T_82 = io_B[4:1]; // @[convert.scala 19:24]
  assign _T_83 = io_B[3:0]; // @[convert.scala 19:43]
  assign _T_84 = _T_82 ^ _T_83; // @[convert.scala 19:39]
  assign _T_85 = _T_84[3:2]; // @[LZD.scala 43:32]
  assign _T_86 = _T_85 != 2'h0; // @[LZD.scala 39:14]
  assign _T_87 = _T_85[1]; // @[LZD.scala 39:21]
  assign _T_88 = _T_85[0]; // @[LZD.scala 39:30]
  assign _T_89 = ~ _T_88; // @[LZD.scala 39:27]
  assign _T_90 = _T_87 | _T_89; // @[LZD.scala 39:25]
  assign _T_91 = {_T_86,_T_90}; // @[Cat.scala 29:58]
  assign _T_92 = _T_84[1:0]; // @[LZD.scala 44:32]
  assign _T_93 = _T_92 != 2'h0; // @[LZD.scala 39:14]
  assign _T_94 = _T_92[1]; // @[LZD.scala 39:21]
  assign _T_95 = _T_92[0]; // @[LZD.scala 39:30]
  assign _T_96 = ~ _T_95; // @[LZD.scala 39:27]
  assign _T_97 = _T_94 | _T_96; // @[LZD.scala 39:25]
  assign _T_98 = {_T_93,_T_97}; // @[Cat.scala 29:58]
  assign _T_99 = _T_91[1]; // @[Shift.scala 12:21]
  assign _T_100 = _T_98[1]; // @[Shift.scala 12:21]
  assign _T_101 = _T_99 | _T_100; // @[LZD.scala 49:16]
  assign _T_102 = ~ _T_100; // @[LZD.scala 49:27]
  assign _T_103 = _T_99 | _T_102; // @[LZD.scala 49:25]
  assign _T_104 = _T_91[0:0]; // @[LZD.scala 49:47]
  assign _T_105 = _T_98[0:0]; // @[LZD.scala 49:59]
  assign _T_106 = _T_99 ? _T_104 : _T_105; // @[LZD.scala 49:35]
  assign _T_108 = {_T_101,_T_103,_T_106}; // @[Cat.scala 29:58]
  assign _T_109 = ~ _T_108; // @[convert.scala 21:22]
  assign _T_110 = io_B[2:0]; // @[convert.scala 22:36]
  assign _T_111 = _T_109 < 3'h3; // @[Shift.scala 16:24]
  assign _T_112 = _T_109[1:0]; // @[Shift.scala 17:37]
  assign _T_113 = _T_112[1]; // @[Shift.scala 12:21]
  assign _T_114 = _T_110[0:0]; // @[Shift.scala 64:52]
  assign _T_116 = {_T_114,2'h0}; // @[Cat.scala 29:58]
  assign _T_117 = _T_113 ? _T_116 : _T_110; // @[Shift.scala 64:27]
  assign _T_118 = _T_112[0:0]; // @[Shift.scala 66:70]
  assign _T_120 = _T_117[1:0]; // @[Shift.scala 64:52]
  assign _T_121 = {_T_120,1'h0}; // @[Cat.scala 29:58]
  assign _T_122 = _T_118 ? _T_121 : _T_117; // @[Shift.scala 64:27]
  assign decB_fraction = _T_111 ? _T_122 : 3'h0; // @[Shift.scala 16:10]
  assign _T_126 = _T_81 == 1'h0; // @[convert.scala 25:26]
  assign _T_128 = _T_81 ? _T_109 : _T_108; // @[convert.scala 25:42]
  assign _T_129 = {_T_126,_T_128}; // @[Cat.scala 29:58]
  assign _T_131 = io_B[4:0]; // @[convert.scala 29:56]
  assign _T_132 = _T_131 != 5'h0; // @[convert.scala 29:60]
  assign _T_133 = ~ _T_132; // @[convert.scala 29:41]
  assign decB_isNaR = _T_79 & _T_133; // @[convert.scala 29:39]
  assign _T_136 = _T_79 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_136 & _T_133; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_129); // @[convert.scala 32:24]
  assign _T_145 = realC[5]; // @[convert.scala 18:24]
  assign _T_146 = realC[4]; // @[convert.scala 18:40]
  assign _T_147 = _T_145 ^ _T_146; // @[convert.scala 18:36]
  assign _T_148 = realC[4:1]; // @[convert.scala 19:24]
  assign _T_149 = realC[3:0]; // @[convert.scala 19:43]
  assign _T_150 = _T_148 ^ _T_149; // @[convert.scala 19:39]
  assign _T_151 = _T_150[3:2]; // @[LZD.scala 43:32]
  assign _T_152 = _T_151 != 2'h0; // @[LZD.scala 39:14]
  assign _T_153 = _T_151[1]; // @[LZD.scala 39:21]
  assign _T_154 = _T_151[0]; // @[LZD.scala 39:30]
  assign _T_155 = ~ _T_154; // @[LZD.scala 39:27]
  assign _T_156 = _T_153 | _T_155; // @[LZD.scala 39:25]
  assign _T_157 = {_T_152,_T_156}; // @[Cat.scala 29:58]
  assign _T_158 = _T_150[1:0]; // @[LZD.scala 44:32]
  assign _T_159 = _T_158 != 2'h0; // @[LZD.scala 39:14]
  assign _T_160 = _T_158[1]; // @[LZD.scala 39:21]
  assign _T_161 = _T_158[0]; // @[LZD.scala 39:30]
  assign _T_162 = ~ _T_161; // @[LZD.scala 39:27]
  assign _T_163 = _T_160 | _T_162; // @[LZD.scala 39:25]
  assign _T_164 = {_T_159,_T_163}; // @[Cat.scala 29:58]
  assign _T_165 = _T_157[1]; // @[Shift.scala 12:21]
  assign _T_166 = _T_164[1]; // @[Shift.scala 12:21]
  assign _T_167 = _T_165 | _T_166; // @[LZD.scala 49:16]
  assign _T_168 = ~ _T_166; // @[LZD.scala 49:27]
  assign _T_169 = _T_165 | _T_168; // @[LZD.scala 49:25]
  assign _T_170 = _T_157[0:0]; // @[LZD.scala 49:47]
  assign _T_171 = _T_164[0:0]; // @[LZD.scala 49:59]
  assign _T_172 = _T_165 ? _T_170 : _T_171; // @[LZD.scala 49:35]
  assign _T_174 = {_T_167,_T_169,_T_172}; // @[Cat.scala 29:58]
  assign _T_175 = ~ _T_174; // @[convert.scala 21:22]
  assign _T_176 = realC[2:0]; // @[convert.scala 22:36]
  assign _T_177 = _T_175 < 3'h3; // @[Shift.scala 16:24]
  assign _T_178 = _T_175[1:0]; // @[Shift.scala 17:37]
  assign _T_179 = _T_178[1]; // @[Shift.scala 12:21]
  assign _T_180 = _T_176[0:0]; // @[Shift.scala 64:52]
  assign _T_182 = {_T_180,2'h0}; // @[Cat.scala 29:58]
  assign _T_183 = _T_179 ? _T_182 : _T_176; // @[Shift.scala 64:27]
  assign _T_184 = _T_178[0:0]; // @[Shift.scala 66:70]
  assign _T_186 = _T_183[1:0]; // @[Shift.scala 64:52]
  assign _T_187 = {_T_186,1'h0}; // @[Cat.scala 29:58]
  assign _T_192 = _T_147 == 1'h0; // @[convert.scala 25:26]
  assign _T_194 = _T_147 ? _T_175 : _T_174; // @[convert.scala 25:42]
  assign _T_195 = {_T_192,_T_194}; // @[Cat.scala 29:58]
  assign _T_197 = realC[4:0]; // @[convert.scala 29:56]
  assign _T_198 = _T_197 != 5'h0; // @[convert.scala 29:60]
  assign _T_199 = ~ _T_198; // @[convert.scala 29:41]
  assign decC_isNaR = _T_145 & _T_199; // @[convert.scala 29:39]
  assign _T_202 = _T_145 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_202 & _T_199; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_195); // @[convert.scala 32:24]
  assign _T_210 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_210 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_211 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_212 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_213 = _T_211 & _T_212; // @[PositFMA.scala 59:45]
  assign _T_215 = {_T_13,_T_213,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_215); // @[PositFMA.scala 59:76]
  assign _T_216 = ~ _T_79; // @[PositFMA.scala 60:34]
  assign _T_217 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_218 = _T_216 & _T_217; // @[PositFMA.scala 60:45]
  assign _T_220 = {_T_79,_T_218,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_220); // @[PositFMA.scala 60:76]
  assign _T_221 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 62:25]
  assign sigP = $unsigned(_T_221); // @[PositFMA.scala 62:33]
  assign head2 = sigP[9:8]; // @[PositFMA.scala 63:28]
  assign _T_222 = head2[1]; // @[PositFMA.scala 64:31]
  assign _T_223 = ~ _T_222; // @[PositFMA.scala 64:25]
  assign _T_224 = head2[0]; // @[PositFMA.scala 64:42]
  assign addTwo = _T_223 & _T_224; // @[PositFMA.scala 64:35]
  assign _T_225 = sigP[9]; // @[PositFMA.scala 66:23]
  assign _T_226 = sigP[7]; // @[PositFMA.scala 66:49]
  assign addOne = _T_225 ^ _T_226; // @[PositFMA.scala 66:43]
  assign _T_227 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_227)}; // @[PositFMA.scala 67:39]
  assign mulSign = sigP[9:9]; // @[PositFMA.scala 68:28]
  assign _T_228 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 70:30]
  assign _GEN_12 = {{2{expBias[2]}},expBias}; // @[PositFMA.scala 70:44]
  assign _T_230 = $signed(_T_228) + $signed(_GEN_12); // @[PositFMA.scala 70:44]
  assign mulScale = $signed(_T_230); // @[PositFMA.scala 70:44]
  assign _T_231 = sigP[7:0]; // @[PositFMA.scala 73:29]
  assign _T_232 = sigP[6:0]; // @[PositFMA.scala 74:29]
  assign _T_233 = {_T_232, 1'h0}; // @[PositFMA.scala 74:48]
  assign mulSigTmp = addOne ? _T_231 : _T_233; // @[PositFMA.scala 71:22]
  assign _T_235 = mulSigTmp[7:7]; // @[PositFMA.scala 78:39]
  assign _T_236 = _T_235 | addTwo; // @[PositFMA.scala 78:43]
  assign _T_237 = mulSigTmp[6:0]; // @[PositFMA.scala 79:39]
  assign mulSig = {mulSign,_T_236,_T_237}; // @[Cat.scala 29:58]
  assign _T_263 = ~ addSign_phase2; // @[PositFMA.scala 108:29]
  assign _T_264 = ~ addZero_phase2; // @[PositFMA.scala 108:47]
  assign _T_265 = _T_263 & _T_264; // @[PositFMA.scala 108:45]
  assign extAddSig = {addSign_phase2,_T_265,addFrac_phase2,4'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[3]}},addScale_phase2}; // @[PositFMA.scala 112:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 112:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[3]}},addScale_phase2}); // @[PositFMA.scala 113:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[3]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 114:26]
  assign _T_269 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 115:36]
  assign scaleDiff = $signed(_T_269); // @[PositFMA.scala 115:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 116:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 117:26]
  assign _T_270 = $unsigned(scaleDiff); // @[PositFMA.scala 118:69]
  assign _T_271 = _T_270 < 5'h9; // @[Shift.scala 39:24]
  assign _T_272 = _T_270[3:0]; // @[Shift.scala 40:44]
  assign _T_273 = smallerSigTmp[8:8]; // @[Shift.scala 90:30]
  assign _T_274 = smallerSigTmp[7:0]; // @[Shift.scala 90:48]
  assign _T_275 = _T_274 != 8'h0; // @[Shift.scala 90:57]
  assign _T_276 = _T_273 | _T_275; // @[Shift.scala 90:39]
  assign _T_277 = _T_272[3]; // @[Shift.scala 12:21]
  assign _T_278 = smallerSigTmp[8]; // @[Shift.scala 12:21]
  assign _T_280 = _T_278 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_281 = {_T_280,_T_276}; // @[Cat.scala 29:58]
  assign _T_282 = _T_277 ? _T_281 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_283 = _T_272[2:0]; // @[Shift.scala 92:77]
  assign _T_284 = _T_282[8:4]; // @[Shift.scala 90:30]
  assign _T_285 = _T_282[3:0]; // @[Shift.scala 90:48]
  assign _T_286 = _T_285 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{4'd0}, _T_286}; // @[Shift.scala 90:39]
  assign _T_287 = _T_284 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_288 = _T_283[2]; // @[Shift.scala 12:21]
  assign _T_289 = _T_282[8]; // @[Shift.scala 12:21]
  assign _T_291 = _T_289 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_292 = {_T_291,_T_287}; // @[Cat.scala 29:58]
  assign _T_293 = _T_288 ? _T_292 : _T_282; // @[Shift.scala 91:22]
  assign _T_294 = _T_283[1:0]; // @[Shift.scala 92:77]
  assign _T_295 = _T_293[8:2]; // @[Shift.scala 90:30]
  assign _T_296 = _T_293[1:0]; // @[Shift.scala 90:48]
  assign _T_297 = _T_296 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{6'd0}, _T_297}; // @[Shift.scala 90:39]
  assign _T_298 = _T_295 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_299 = _T_294[1]; // @[Shift.scala 12:21]
  assign _T_300 = _T_293[8]; // @[Shift.scala 12:21]
  assign _T_302 = _T_300 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_303 = {_T_302,_T_298}; // @[Cat.scala 29:58]
  assign _T_304 = _T_299 ? _T_303 : _T_293; // @[Shift.scala 91:22]
  assign _T_305 = _T_294[0:0]; // @[Shift.scala 92:77]
  assign _T_306 = _T_304[8:1]; // @[Shift.scala 90:30]
  assign _T_307 = _T_304[0:0]; // @[Shift.scala 90:48]
  assign _GEN_16 = {{7'd0}, _T_307}; // @[Shift.scala 90:39]
  assign _T_309 = _T_306 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_311 = _T_304[8]; // @[Shift.scala 12:21]
  assign _T_312 = {_T_311,_T_309}; // @[Cat.scala 29:58]
  assign _T_313 = _T_305 ? _T_312 : _T_304; // @[Shift.scala 91:22]
  assign _T_316 = _T_278 ? 9'h1ff : 9'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_271 ? _T_313 : _T_316; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 119:34]
  assign _T_317 = mulSig_phase2[8:8]; // @[PositFMA.scala 120:42]
  assign _T_318 = _T_317 ^ addSign_phase2; // @[PositFMA.scala 120:46]
  assign _T_319 = rawSumSig[9:9]; // @[PositFMA.scala 120:79]
  assign sumSign = _T_318 ^ _T_319; // @[PositFMA.scala 120:63]
  assign _T_321 = greaterSig + smallerSig; // @[PositFMA.scala 121:50]
  assign signSumSig = {sumSign,_T_321}; // @[Cat.scala 29:58]
  assign _T_322 = signSumSig[9:1]; // @[PositFMA.scala 126:33]
  assign _T_323 = signSumSig[8:0]; // @[PositFMA.scala 126:68]
  assign sumXor = _T_322 ^ _T_323; // @[PositFMA.scala 126:51]
  assign _T_324 = sumXor[8:1]; // @[LZD.scala 43:32]
  assign _T_325 = _T_324[7:4]; // @[LZD.scala 43:32]
  assign _T_326 = _T_325[3:2]; // @[LZD.scala 43:32]
  assign _T_327 = _T_326 != 2'h0; // @[LZD.scala 39:14]
  assign _T_328 = _T_326[1]; // @[LZD.scala 39:21]
  assign _T_329 = _T_326[0]; // @[LZD.scala 39:30]
  assign _T_330 = ~ _T_329; // @[LZD.scala 39:27]
  assign _T_331 = _T_328 | _T_330; // @[LZD.scala 39:25]
  assign _T_332 = {_T_327,_T_331}; // @[Cat.scala 29:58]
  assign _T_333 = _T_325[1:0]; // @[LZD.scala 44:32]
  assign _T_334 = _T_333 != 2'h0; // @[LZD.scala 39:14]
  assign _T_335 = _T_333[1]; // @[LZD.scala 39:21]
  assign _T_336 = _T_333[0]; // @[LZD.scala 39:30]
  assign _T_337 = ~ _T_336; // @[LZD.scala 39:27]
  assign _T_338 = _T_335 | _T_337; // @[LZD.scala 39:25]
  assign _T_339 = {_T_334,_T_338}; // @[Cat.scala 29:58]
  assign _T_340 = _T_332[1]; // @[Shift.scala 12:21]
  assign _T_341 = _T_339[1]; // @[Shift.scala 12:21]
  assign _T_342 = _T_340 | _T_341; // @[LZD.scala 49:16]
  assign _T_343 = ~ _T_341; // @[LZD.scala 49:27]
  assign _T_344 = _T_340 | _T_343; // @[LZD.scala 49:25]
  assign _T_345 = _T_332[0:0]; // @[LZD.scala 49:47]
  assign _T_346 = _T_339[0:0]; // @[LZD.scala 49:59]
  assign _T_347 = _T_340 ? _T_345 : _T_346; // @[LZD.scala 49:35]
  assign _T_349 = {_T_342,_T_344,_T_347}; // @[Cat.scala 29:58]
  assign _T_350 = _T_324[3:0]; // @[LZD.scala 44:32]
  assign _T_351 = _T_350[3:2]; // @[LZD.scala 43:32]
  assign _T_352 = _T_351 != 2'h0; // @[LZD.scala 39:14]
  assign _T_353 = _T_351[1]; // @[LZD.scala 39:21]
  assign _T_354 = _T_351[0]; // @[LZD.scala 39:30]
  assign _T_355 = ~ _T_354; // @[LZD.scala 39:27]
  assign _T_356 = _T_353 | _T_355; // @[LZD.scala 39:25]
  assign _T_357 = {_T_352,_T_356}; // @[Cat.scala 29:58]
  assign _T_358 = _T_350[1:0]; // @[LZD.scala 44:32]
  assign _T_359 = _T_358 != 2'h0; // @[LZD.scala 39:14]
  assign _T_360 = _T_358[1]; // @[LZD.scala 39:21]
  assign _T_361 = _T_358[0]; // @[LZD.scala 39:30]
  assign _T_362 = ~ _T_361; // @[LZD.scala 39:27]
  assign _T_363 = _T_360 | _T_362; // @[LZD.scala 39:25]
  assign _T_364 = {_T_359,_T_363}; // @[Cat.scala 29:58]
  assign _T_365 = _T_357[1]; // @[Shift.scala 12:21]
  assign _T_366 = _T_364[1]; // @[Shift.scala 12:21]
  assign _T_367 = _T_365 | _T_366; // @[LZD.scala 49:16]
  assign _T_368 = ~ _T_366; // @[LZD.scala 49:27]
  assign _T_369 = _T_365 | _T_368; // @[LZD.scala 49:25]
  assign _T_370 = _T_357[0:0]; // @[LZD.scala 49:47]
  assign _T_371 = _T_364[0:0]; // @[LZD.scala 49:59]
  assign _T_372 = _T_365 ? _T_370 : _T_371; // @[LZD.scala 49:35]
  assign _T_374 = {_T_367,_T_369,_T_372}; // @[Cat.scala 29:58]
  assign _T_375 = _T_349[2]; // @[Shift.scala 12:21]
  assign _T_376 = _T_374[2]; // @[Shift.scala 12:21]
  assign _T_377 = _T_375 | _T_376; // @[LZD.scala 49:16]
  assign _T_378 = ~ _T_376; // @[LZD.scala 49:27]
  assign _T_379 = _T_375 | _T_378; // @[LZD.scala 49:25]
  assign _T_380 = _T_349[1:0]; // @[LZD.scala 49:47]
  assign _T_381 = _T_374[1:0]; // @[LZD.scala 49:59]
  assign _T_382 = _T_375 ? _T_380 : _T_381; // @[LZD.scala 49:35]
  assign _T_384 = {_T_377,_T_379,_T_382}; // @[Cat.scala 29:58]
  assign _T_385 = sumXor[0:0]; // @[LZD.scala 44:32]
  assign _T_387 = _T_384[3]; // @[Shift.scala 12:21]
  assign _T_390 = {2'h3,_T_385}; // @[Cat.scala 29:58]
  assign _T_391 = _T_384[2:0]; // @[LZD.scala 55:32]
  assign _T_392 = _T_387 ? _T_391 : _T_390; // @[LZD.scala 55:20]
  assign sumLZD = {_T_387,_T_392}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 128:24]
  assign _T_393 = signSumSig[7:0]; // @[PositFMA.scala 129:38]
  assign _T_394 = shiftValue < 4'h8; // @[Shift.scala 16:24]
  assign _T_395 = shiftValue[2:0]; // @[Shift.scala 17:37]
  assign _T_396 = _T_395[2]; // @[Shift.scala 12:21]
  assign _T_397 = _T_393[3:0]; // @[Shift.scala 64:52]
  assign _T_399 = {_T_397,4'h0}; // @[Cat.scala 29:58]
  assign _T_400 = _T_396 ? _T_399 : _T_393; // @[Shift.scala 64:27]
  assign _T_401 = _T_395[1:0]; // @[Shift.scala 66:70]
  assign _T_402 = _T_401[1]; // @[Shift.scala 12:21]
  assign _T_403 = _T_400[5:0]; // @[Shift.scala 64:52]
  assign _T_405 = {_T_403,2'h0}; // @[Cat.scala 29:58]
  assign _T_406 = _T_402 ? _T_405 : _T_400; // @[Shift.scala 64:27]
  assign _T_407 = _T_401[0:0]; // @[Shift.scala 66:70]
  assign _T_409 = _T_406[6:0]; // @[Shift.scala 64:52]
  assign _T_410 = {_T_409,1'h0}; // @[Cat.scala 29:58]
  assign _T_411 = _T_407 ? _T_410 : _T_406; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_394 ? _T_411 : 8'h0; // @[Shift.scala 16:10]
  assign _T_413 = $signed(greaterScale) + $signed(5'sh2); // @[PositFMA.scala 132:36]
  assign _T_414 = $signed(_T_413); // @[PositFMA.scala 132:36]
  assign _T_415 = {1'h1,_T_387,_T_392}; // @[Cat.scala 29:58]
  assign _T_416 = $signed(_T_415); // @[PositFMA.scala 132:61]
  assign _T_418 = $signed(_T_414) + $signed(_T_416); // @[PositFMA.scala 132:42]
  assign sumScale = $signed(_T_418); // @[PositFMA.scala 132:42]
  assign sumFrac = normalFracTmp[7:5]; // @[PositFMA.scala 133:41]
  assign grsTmp = normalFracTmp[4:0]; // @[PositFMA.scala 136:41]
  assign _T_419 = grsTmp[4:3]; // @[PositFMA.scala 139:40]
  assign _T_420 = grsTmp[2:0]; // @[PositFMA.scala 139:56]
  assign _T_421 = _T_420 != 3'h0; // @[PositFMA.scala 139:60]
  assign underflow = $signed(sumScale) < $signed(-5'sh5); // @[PositFMA.scala 146:32]
  assign overflow = $signed(sumScale) > $signed(5'sh4); // @[PositFMA.scala 147:32]
  assign _T_422 = signSumSig != 10'h0; // @[PositFMA.scala 156:32]
  assign decF_isZero = ~ _T_422; // @[PositFMA.scala 156:20]
  assign _T_424 = underflow ? $signed(-5'sh5) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_425 = overflow ? $signed(5'sh4) : $signed(_T_424); // @[Mux.scala 87:16]
  assign _GEN_17 = _T_425[3:0]; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  assign decF_scale = $signed(_GEN_17); // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  assign _T_427 = decF_scale[3:3]; // @[convert.scala 49:36]
  assign _T_429 = ~ decF_scale; // @[convert.scala 50:36]
  assign _T_430 = $signed(_T_429); // @[convert.scala 50:36]
  assign _T_431 = _T_427 ? $signed(_T_430) : $signed(decF_scale); // @[convert.scala 50:28]
  assign _T_432 = _T_427 ^ sumSign; // @[convert.scala 51:31]
  assign _T_433 = ~ _T_432; // @[convert.scala 53:34]
  assign _T_436 = {_T_433,_T_432,sumFrac,_T_419,_T_421}; // @[Cat.scala 29:58]
  assign _T_437 = $unsigned(_T_431); // @[Shift.scala 39:17]
  assign _T_438 = _T_437 < 4'h8; // @[Shift.scala 39:24]
  assign _T_439 = _T_431[2:0]; // @[Shift.scala 40:44]
  assign _T_440 = _T_436[7:4]; // @[Shift.scala 90:30]
  assign _T_441 = _T_436[3:0]; // @[Shift.scala 90:48]
  assign _T_442 = _T_441 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_18 = {{3'd0}, _T_442}; // @[Shift.scala 90:39]
  assign _T_443 = _T_440 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_444 = _T_439[2]; // @[Shift.scala 12:21]
  assign _T_445 = _T_436[7]; // @[Shift.scala 12:21]
  assign _T_447 = _T_445 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_448 = {_T_447,_T_443}; // @[Cat.scala 29:58]
  assign _T_449 = _T_444 ? _T_448 : _T_436; // @[Shift.scala 91:22]
  assign _T_450 = _T_439[1:0]; // @[Shift.scala 92:77]
  assign _T_451 = _T_449[7:2]; // @[Shift.scala 90:30]
  assign _T_452 = _T_449[1:0]; // @[Shift.scala 90:48]
  assign _T_453 = _T_452 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_19 = {{5'd0}, _T_453}; // @[Shift.scala 90:39]
  assign _T_454 = _T_451 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_455 = _T_450[1]; // @[Shift.scala 12:21]
  assign _T_456 = _T_449[7]; // @[Shift.scala 12:21]
  assign _T_458 = _T_456 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_459 = {_T_458,_T_454}; // @[Cat.scala 29:58]
  assign _T_460 = _T_455 ? _T_459 : _T_449; // @[Shift.scala 91:22]
  assign _T_461 = _T_450[0:0]; // @[Shift.scala 92:77]
  assign _T_462 = _T_460[7:1]; // @[Shift.scala 90:30]
  assign _T_463 = _T_460[0:0]; // @[Shift.scala 90:48]
  assign _GEN_20 = {{6'd0}, _T_463}; // @[Shift.scala 90:39]
  assign _T_465 = _T_462 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_467 = _T_460[7]; // @[Shift.scala 12:21]
  assign _T_468 = {_T_467,_T_465}; // @[Cat.scala 29:58]
  assign _T_469 = _T_461 ? _T_468 : _T_460; // @[Shift.scala 91:22]
  assign _T_472 = _T_445 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_473 = _T_438 ? _T_469 : _T_472; // @[Shift.scala 39:10]
  assign _T_474 = _T_473[3]; // @[convert.scala 55:31]
  assign _T_475 = _T_473[2]; // @[convert.scala 56:31]
  assign _T_476 = _T_473[1]; // @[convert.scala 57:31]
  assign _T_477 = _T_473[0]; // @[convert.scala 58:31]
  assign _T_478 = _T_473[7:3]; // @[convert.scala 59:69]
  assign _T_479 = _T_478 != 5'h0; // @[convert.scala 59:81]
  assign _T_480 = ~ _T_479; // @[convert.scala 59:50]
  assign _T_482 = _T_478 == 5'h1f; // @[convert.scala 60:81]
  assign _T_483 = _T_474 | _T_476; // @[convert.scala 61:44]
  assign _T_484 = _T_483 | _T_477; // @[convert.scala 61:52]
  assign _T_485 = _T_475 & _T_484; // @[convert.scala 61:36]
  assign _T_486 = ~ _T_482; // @[convert.scala 62:63]
  assign _T_487 = _T_486 & _T_485; // @[convert.scala 62:103]
  assign _T_488 = _T_480 | _T_487; // @[convert.scala 62:60]
  assign _GEN_21 = {{4'd0}, _T_488}; // @[convert.scala 63:56]
  assign _T_491 = _T_478 + _GEN_21; // @[convert.scala 63:56]
  assign _T_492 = {sumSign,_T_491}; // @[Cat.scala 29:58]
  assign io_F = _T_500; // @[PositFMA.scala 176:15]
  assign io_outValid = _T_496; // @[PositFMA.scala 175:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulSig_phase2 = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_496 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_500 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      if (_T_177) begin
        if (_T_184) begin
          addFrac_phase2 <= _T_187;
        end else begin
          if (_T_179) begin
            addFrac_phase2 <= _T_182;
          end else begin
            addFrac_phase2 <= _T_176;
          end
        end
      end else begin
        addFrac_phase2 <= 3'h0;
      end
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_145;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_496 <= 1'h0;
    end else begin
      _T_496 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_500 <= 6'h20;
      end else begin
        if (decF_isZero) begin
          _T_500 <= 6'h0;
        end else begin
          _T_500 <= _T_492;
        end
      end
    end
  end
endmodule
