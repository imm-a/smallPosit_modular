module Sig_op_approx5_0(
  input        clock,
  input        reset,
  input  [4:0] io_A,
  input  [4:0] io_B,
  output       io_greaterSign,
  output       io_smallerSign,
  output [2:0] io_greaterExp,
  output [3:0] io_greaterSig,
  output [6:0] io_smallerSig,
  output       io_AisNar,
  output       io_BisNar,
  output       io_AisZero,
  output       io_BisZero
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [2:0] _T_4; // @[convert.scala 19:24]
  wire [2:0] _T_5; // @[convert.scala 19:43]
  wire [2:0] _T_6; // @[convert.scala 19:39]
  wire [1:0] _T_7; // @[LZD.scala 43:32]
  wire  _T_8; // @[LZD.scala 39:14]
  wire  _T_9; // @[LZD.scala 39:21]
  wire  _T_10; // @[LZD.scala 39:30]
  wire  _T_11; // @[LZD.scala 39:27]
  wire  _T_12; // @[LZD.scala 39:25]
  wire [1:0] _T_13; // @[Cat.scala 29:58]
  wire  _T_14; // @[LZD.scala 44:32]
  wire  _T_16; // @[Shift.scala 12:21]
  wire  _T_18; // @[LZD.scala 55:32]
  wire  _T_19; // @[LZD.scala 55:20]
  wire [1:0] _T_20; // @[Cat.scala 29:58]
  wire [1:0] _T_21; // @[convert.scala 21:22]
  wire [1:0] _T_22; // @[convert.scala 22:36]
  wire  _T_23; // @[Shift.scala 16:24]
  wire  _T_24; // @[Shift.scala 17:37]
  wire  _T_26; // @[Shift.scala 64:52]
  wire [1:0] _T_27; // @[Cat.scala 29:58]
  wire [1:0] _T_28; // @[Shift.scala 64:27]
  wire [1:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_32; // @[convert.scala 25:26]
  wire [1:0] _T_34; // @[convert.scala 25:42]
  wire [2:0] _T_35; // @[Cat.scala 29:58]
  wire [3:0] _T_37; // @[convert.scala 29:56]
  wire  _T_38; // @[convert.scala 29:60]
  wire  _T_39; // @[convert.scala 29:41]
  wire  _T_42; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [2:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_51; // @[convert.scala 18:24]
  wire  _T_52; // @[convert.scala 18:40]
  wire  _T_53; // @[convert.scala 18:36]
  wire [2:0] _T_54; // @[convert.scala 19:24]
  wire [2:0] _T_55; // @[convert.scala 19:43]
  wire [2:0] _T_56; // @[convert.scala 19:39]
  wire [1:0] _T_57; // @[LZD.scala 43:32]
  wire  _T_58; // @[LZD.scala 39:14]
  wire  _T_59; // @[LZD.scala 39:21]
  wire  _T_60; // @[LZD.scala 39:30]
  wire  _T_61; // @[LZD.scala 39:27]
  wire  _T_62; // @[LZD.scala 39:25]
  wire [1:0] _T_63; // @[Cat.scala 29:58]
  wire  _T_64; // @[LZD.scala 44:32]
  wire  _T_66; // @[Shift.scala 12:21]
  wire  _T_68; // @[LZD.scala 55:32]
  wire  _T_69; // @[LZD.scala 55:20]
  wire [1:0] _T_70; // @[Cat.scala 29:58]
  wire [1:0] _T_71; // @[convert.scala 21:22]
  wire [1:0] _T_72; // @[convert.scala 22:36]
  wire  _T_73; // @[Shift.scala 16:24]
  wire  _T_74; // @[Shift.scala 17:37]
  wire  _T_76; // @[Shift.scala 64:52]
  wire [1:0] _T_77; // @[Cat.scala 29:58]
  wire [1:0] _T_78; // @[Shift.scala 64:27]
  wire [1:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_82; // @[convert.scala 25:26]
  wire [1:0] _T_84; // @[convert.scala 25:42]
  wire [2:0] _T_85; // @[Cat.scala 29:58]
  wire [3:0] _T_87; // @[convert.scala 29:56]
  wire  _T_88; // @[convert.scala 29:60]
  wire  _T_89; // @[convert.scala 29:41]
  wire  _T_92; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [2:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_101; // @[Sig_op_approx.scala 37:30]
  wire [2:0] scale_diff; // @[Sig_op_approx.scala 37:30]
  wire  _T_102; // @[Sig_op_approx.scala 38:37]
  wire  aGTb; // @[Sig_op_approx.scala 38:21]
  wire [1:0] greaterFrac; // @[Sig_op_approx.scala 43:24]
  wire [1:0] smallerFrac; // @[Sig_op_approx.scala 44:24]
  wire  smallerZero; // @[Sig_op_approx.scala 45:24]
  wire [2:0] _T_108; // @[Sig_op_approx.scala 46:35]
  wire [2:0] _T_109; // @[Sig_op_approx.scala 46:35]
  wire [2:0] sdiff; // @[Sig_op_approx.scala 46:18]
  wire  _T_110; // @[Sig_op_approx.scala 51:53]
  wire  _T_111; // @[Sig_op_approx.scala 51:36]
  wire [6:0] _T_114; // @[Cat.scala 29:58]
  wire [2:0] _T_115; // @[Sig_op_approx.scala 51:119]
  wire  _T_116; // @[Shift.scala 39:24]
  wire [2:0] _T_118; // @[Shift.scala 90:30]
  wire [3:0] _T_119; // @[Shift.scala 90:48]
  wire  _T_120; // @[Shift.scala 90:57]
  wire [2:0] _GEN_0; // @[Shift.scala 90:39]
  wire [2:0] _T_121; // @[Shift.scala 90:39]
  wire  _T_122; // @[Shift.scala 12:21]
  wire  _T_123; // @[Shift.scala 12:21]
  wire [3:0] _T_125; // @[Bitwise.scala 71:12]
  wire [6:0] _T_126; // @[Cat.scala 29:58]
  wire [6:0] _T_127; // @[Shift.scala 91:22]
  wire [1:0] _T_128; // @[Shift.scala 92:77]
  wire [4:0] _T_129; // @[Shift.scala 90:30]
  wire [1:0] _T_130; // @[Shift.scala 90:48]
  wire  _T_131; // @[Shift.scala 90:57]
  wire [4:0] _GEN_1; // @[Shift.scala 90:39]
  wire [4:0] _T_132; // @[Shift.scala 90:39]
  wire  _T_133; // @[Shift.scala 12:21]
  wire  _T_134; // @[Shift.scala 12:21]
  wire [1:0] _T_136; // @[Bitwise.scala 71:12]
  wire [6:0] _T_137; // @[Cat.scala 29:58]
  wire [6:0] _T_138; // @[Shift.scala 91:22]
  wire  _T_139; // @[Shift.scala 92:77]
  wire [5:0] _T_140; // @[Shift.scala 90:30]
  wire  _T_141; // @[Shift.scala 90:48]
  wire [5:0] _GEN_2; // @[Shift.scala 90:39]
  wire [5:0] _T_143; // @[Shift.scala 90:39]
  wire  _T_145; // @[Shift.scala 12:21]
  wire [6:0] _T_146; // @[Cat.scala 29:58]
  wire [6:0] _T_147; // @[Shift.scala 91:22]
  wire [6:0] _T_150; // @[Bitwise.scala 71:12]
  wire  _T_151; // @[Sig_op_approx.scala 57:40]
  wire [1:0] _T_152; // @[Cat.scala 29:58]
  assign _T_1 = io_A[4]; // @[convert.scala 18:24]
  assign _T_2 = io_A[3]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[3:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[2:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[2:1]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7 != 2'h0; // @[LZD.scala 39:14]
  assign _T_9 = _T_7[1]; // @[LZD.scala 39:21]
  assign _T_10 = _T_7[0]; // @[LZD.scala 39:30]
  assign _T_11 = ~ _T_10; // @[LZD.scala 39:27]
  assign _T_12 = _T_9 | _T_11; // @[LZD.scala 39:25]
  assign _T_13 = {_T_8,_T_12}; // @[Cat.scala 29:58]
  assign _T_14 = _T_6[0:0]; // @[LZD.scala 44:32]
  assign _T_16 = _T_13[1]; // @[Shift.scala 12:21]
  assign _T_18 = _T_13[0:0]; // @[LZD.scala 55:32]
  assign _T_19 = _T_16 ? _T_18 : _T_14; // @[LZD.scala 55:20]
  assign _T_20 = {_T_16,_T_19}; // @[Cat.scala 29:58]
  assign _T_21 = ~ _T_20; // @[convert.scala 21:22]
  assign _T_22 = io_A[1:0]; // @[convert.scala 22:36]
  assign _T_23 = _T_21 < 2'h2; // @[Shift.scala 16:24]
  assign _T_24 = _T_21[0]; // @[Shift.scala 17:37]
  assign _T_26 = _T_22[0:0]; // @[Shift.scala 64:52]
  assign _T_27 = {_T_26,1'h0}; // @[Cat.scala 29:58]
  assign _T_28 = _T_24 ? _T_27 : _T_22; // @[Shift.scala 64:27]
  assign decA_fraction = _T_23 ? _T_28 : 2'h0; // @[Shift.scala 16:10]
  assign _T_32 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_34 = _T_3 ? _T_21 : _T_20; // @[convert.scala 25:42]
  assign _T_35 = {_T_32,_T_34}; // @[Cat.scala 29:58]
  assign _T_37 = io_A[3:0]; // @[convert.scala 29:56]
  assign _T_38 = _T_37 != 4'h0; // @[convert.scala 29:60]
  assign _T_39 = ~ _T_38; // @[convert.scala 29:41]
  assign _T_42 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_42 & _T_39; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_35); // @[convert.scala 32:24]
  assign _T_51 = io_B[4]; // @[convert.scala 18:24]
  assign _T_52 = io_B[3]; // @[convert.scala 18:40]
  assign _T_53 = _T_51 ^ _T_52; // @[convert.scala 18:36]
  assign _T_54 = io_B[3:1]; // @[convert.scala 19:24]
  assign _T_55 = io_B[2:0]; // @[convert.scala 19:43]
  assign _T_56 = _T_54 ^ _T_55; // @[convert.scala 19:39]
  assign _T_57 = _T_56[2:1]; // @[LZD.scala 43:32]
  assign _T_58 = _T_57 != 2'h0; // @[LZD.scala 39:14]
  assign _T_59 = _T_57[1]; // @[LZD.scala 39:21]
  assign _T_60 = _T_57[0]; // @[LZD.scala 39:30]
  assign _T_61 = ~ _T_60; // @[LZD.scala 39:27]
  assign _T_62 = _T_59 | _T_61; // @[LZD.scala 39:25]
  assign _T_63 = {_T_58,_T_62}; // @[Cat.scala 29:58]
  assign _T_64 = _T_56[0:0]; // @[LZD.scala 44:32]
  assign _T_66 = _T_63[1]; // @[Shift.scala 12:21]
  assign _T_68 = _T_63[0:0]; // @[LZD.scala 55:32]
  assign _T_69 = _T_66 ? _T_68 : _T_64; // @[LZD.scala 55:20]
  assign _T_70 = {_T_66,_T_69}; // @[Cat.scala 29:58]
  assign _T_71 = ~ _T_70; // @[convert.scala 21:22]
  assign _T_72 = io_B[1:0]; // @[convert.scala 22:36]
  assign _T_73 = _T_71 < 2'h2; // @[Shift.scala 16:24]
  assign _T_74 = _T_71[0]; // @[Shift.scala 17:37]
  assign _T_76 = _T_72[0:0]; // @[Shift.scala 64:52]
  assign _T_77 = {_T_76,1'h0}; // @[Cat.scala 29:58]
  assign _T_78 = _T_74 ? _T_77 : _T_72; // @[Shift.scala 64:27]
  assign decB_fraction = _T_73 ? _T_78 : 2'h0; // @[Shift.scala 16:10]
  assign _T_82 = _T_53 == 1'h0; // @[convert.scala 25:26]
  assign _T_84 = _T_53 ? _T_71 : _T_70; // @[convert.scala 25:42]
  assign _T_85 = {_T_82,_T_84}; // @[Cat.scala 29:58]
  assign _T_87 = io_B[3:0]; // @[convert.scala 29:56]
  assign _T_88 = _T_87 != 4'h0; // @[convert.scala 29:60]
  assign _T_89 = ~ _T_88; // @[convert.scala 29:41]
  assign _T_92 = _T_51 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_92 & _T_89; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_85); // @[convert.scala 32:24]
  assign _T_101 = $signed(decA_scale) - $signed(decB_scale); // @[Sig_op_approx.scala 37:30]
  assign scale_diff = $signed(_T_101); // @[Sig_op_approx.scala 37:30]
  assign _T_102 = scale_diff[2:2]; // @[Sig_op_approx.scala 38:37]
  assign aGTb = ~ _T_102; // @[Sig_op_approx.scala 38:21]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[Sig_op_approx.scala 43:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[Sig_op_approx.scala 44:24]
  assign smallerZero = aGTb ? decB_isZero : decA_isZero; // @[Sig_op_approx.scala 45:24]
  assign _T_108 = $signed(3'sh0) - $signed(scale_diff); // @[Sig_op_approx.scala 46:35]
  assign _T_109 = $signed(_T_108); // @[Sig_op_approx.scala 46:35]
  assign sdiff = aGTb ? $signed(scale_diff) : $signed(_T_109); // @[Sig_op_approx.scala 46:18]
  assign _T_110 = io_smallerSign | smallerZero; // @[Sig_op_approx.scala 51:53]
  assign _T_111 = ~ _T_110; // @[Sig_op_approx.scala 51:36]
  assign _T_114 = {io_smallerSign,_T_111,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_115 = $unsigned(sdiff); // @[Sig_op_approx.scala 51:119]
  assign _T_116 = _T_115 < 3'h7; // @[Shift.scala 39:24]
  assign _T_118 = _T_114[6:4]; // @[Shift.scala 90:30]
  assign _T_119 = _T_114[3:0]; // @[Shift.scala 90:48]
  assign _T_120 = _T_119 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{2'd0}, _T_120}; // @[Shift.scala 90:39]
  assign _T_121 = _T_118 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_122 = _T_115[2]; // @[Shift.scala 12:21]
  assign _T_123 = _T_114[6]; // @[Shift.scala 12:21]
  assign _T_125 = _T_123 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_126 = {_T_125,_T_121}; // @[Cat.scala 29:58]
  assign _T_127 = _T_122 ? _T_126 : _T_114; // @[Shift.scala 91:22]
  assign _T_128 = _T_115[1:0]; // @[Shift.scala 92:77]
  assign _T_129 = _T_127[6:2]; // @[Shift.scala 90:30]
  assign _T_130 = _T_127[1:0]; // @[Shift.scala 90:48]
  assign _T_131 = _T_130 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{4'd0}, _T_131}; // @[Shift.scala 90:39]
  assign _T_132 = _T_129 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_133 = _T_128[1]; // @[Shift.scala 12:21]
  assign _T_134 = _T_127[6]; // @[Shift.scala 12:21]
  assign _T_136 = _T_134 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_137 = {_T_136,_T_132}; // @[Cat.scala 29:58]
  assign _T_138 = _T_133 ? _T_137 : _T_127; // @[Shift.scala 91:22]
  assign _T_139 = _T_128[0:0]; // @[Shift.scala 92:77]
  assign _T_140 = _T_138[6:1]; // @[Shift.scala 90:30]
  assign _T_141 = _T_138[0:0]; // @[Shift.scala 90:48]
  assign _GEN_2 = {{5'd0}, _T_141}; // @[Shift.scala 90:39]
  assign _T_143 = _T_140 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_145 = _T_138[6]; // @[Shift.scala 12:21]
  assign _T_146 = {_T_145,_T_143}; // @[Cat.scala 29:58]
  assign _T_147 = _T_139 ? _T_146 : _T_138; // @[Shift.scala 91:22]
  assign _T_150 = _T_123 ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign _T_151 = ~ io_greaterSign; // @[Sig_op_approx.scala 57:40]
  assign _T_152 = {io_greaterSign,_T_151}; // @[Cat.scala 29:58]
  assign io_greaterSign = aGTb ? _T_1 : _T_51; // @[Sig_op_approx.scala 39:18]
  assign io_smallerSign = aGTb ? _T_51 : _T_1; // @[Sig_op_approx.scala 40:18]
  assign io_greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[Sig_op_approx.scala 41:18]
  assign io_greaterSig = {_T_152,greaterFrac}; // @[Sig_op_approx.scala 57:17]
  assign io_smallerSig = _T_116 ? _T_147 : _T_150; // @[Sig_op_approx.scala 52:17]
  assign io_AisNar = _T_1 & _T_39; // @[Sig_op_approx.scala 47:13]
  assign io_BisNar = _T_51 & _T_89; // @[Sig_op_approx.scala 48:13]
  assign io_AisZero = _T_42 & _T_39; // @[Sig_op_approx.scala 49:14]
  assign io_BisZero = _T_92 & _T_89; // @[Sig_op_approx.scala 50:14]
endmodule
