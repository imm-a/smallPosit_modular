module FMAEnc8_0(
  input         clock,
  input         reset,
  input         io_inValid_phase2,
  input  [13:0] io_signSumSig,
  input         io_sumSign,
  input  [3:0]  io_greaterScale,
  input         io_outIsNaR_phase2,
  output [7:0]  io_F,
  output        io_outValid
);
  wire [12:0] _T; // @[FMAEnc.scala 35:36]
  wire [12:0] _T_1; // @[FMAEnc.scala 35:74]
  wire [12:0] sumXor; // @[FMAEnc.scala 35:54]
  wire [7:0] _T_2; // @[LZD.scala 43:32]
  wire [3:0] _T_3; // @[LZD.scala 43:32]
  wire [1:0] _T_4; // @[LZD.scala 43:32]
  wire  _T_5; // @[LZD.scala 39:14]
  wire  _T_6; // @[LZD.scala 39:21]
  wire  _T_7; // @[LZD.scala 39:30]
  wire  _T_8; // @[LZD.scala 39:27]
  wire  _T_9; // @[LZD.scala 39:25]
  wire [1:0] _T_10; // @[Cat.scala 29:58]
  wire [1:0] _T_11; // @[LZD.scala 44:32]
  wire  _T_12; // @[LZD.scala 39:14]
  wire  _T_13; // @[LZD.scala 39:21]
  wire  _T_14; // @[LZD.scala 39:30]
  wire  _T_15; // @[LZD.scala 39:27]
  wire  _T_16; // @[LZD.scala 39:25]
  wire [1:0] _T_17; // @[Cat.scala 29:58]
  wire  _T_18; // @[Shift.scala 12:21]
  wire  _T_19; // @[Shift.scala 12:21]
  wire  _T_20; // @[LZD.scala 49:16]
  wire  _T_21; // @[LZD.scala 49:27]
  wire  _T_22; // @[LZD.scala 49:25]
  wire  _T_23; // @[LZD.scala 49:47]
  wire  _T_24; // @[LZD.scala 49:59]
  wire  _T_25; // @[LZD.scala 49:35]
  wire [2:0] _T_27; // @[Cat.scala 29:58]
  wire [3:0] _T_28; // @[LZD.scala 44:32]
  wire [1:0] _T_29; // @[LZD.scala 43:32]
  wire  _T_30; // @[LZD.scala 39:14]
  wire  _T_31; // @[LZD.scala 39:21]
  wire  _T_32; // @[LZD.scala 39:30]
  wire  _T_33; // @[LZD.scala 39:27]
  wire  _T_34; // @[LZD.scala 39:25]
  wire [1:0] _T_35; // @[Cat.scala 29:58]
  wire [1:0] _T_36; // @[LZD.scala 44:32]
  wire  _T_37; // @[LZD.scala 39:14]
  wire  _T_38; // @[LZD.scala 39:21]
  wire  _T_39; // @[LZD.scala 39:30]
  wire  _T_40; // @[LZD.scala 39:27]
  wire  _T_41; // @[LZD.scala 39:25]
  wire [1:0] _T_42; // @[Cat.scala 29:58]
  wire  _T_43; // @[Shift.scala 12:21]
  wire  _T_44; // @[Shift.scala 12:21]
  wire  _T_45; // @[LZD.scala 49:16]
  wire  _T_46; // @[LZD.scala 49:27]
  wire  _T_47; // @[LZD.scala 49:25]
  wire  _T_48; // @[LZD.scala 49:47]
  wire  _T_49; // @[LZD.scala 49:59]
  wire  _T_50; // @[LZD.scala 49:35]
  wire [2:0] _T_52; // @[Cat.scala 29:58]
  wire  _T_53; // @[Shift.scala 12:21]
  wire  _T_54; // @[Shift.scala 12:21]
  wire  _T_55; // @[LZD.scala 49:16]
  wire  _T_56; // @[LZD.scala 49:27]
  wire  _T_57; // @[LZD.scala 49:25]
  wire [1:0] _T_58; // @[LZD.scala 49:47]
  wire [1:0] _T_59; // @[LZD.scala 49:59]
  wire [1:0] _T_60; // @[LZD.scala 49:35]
  wire [3:0] _T_62; // @[Cat.scala 29:58]
  wire [4:0] _T_63; // @[LZD.scala 44:32]
  wire [3:0] _T_64; // @[LZD.scala 43:32]
  wire [1:0] _T_65; // @[LZD.scala 43:32]
  wire  _T_66; // @[LZD.scala 39:14]
  wire  _T_67; // @[LZD.scala 39:21]
  wire  _T_68; // @[LZD.scala 39:30]
  wire  _T_69; // @[LZD.scala 39:27]
  wire  _T_70; // @[LZD.scala 39:25]
  wire [1:0] _T_71; // @[Cat.scala 29:58]
  wire [1:0] _T_72; // @[LZD.scala 44:32]
  wire  _T_73; // @[LZD.scala 39:14]
  wire  _T_74; // @[LZD.scala 39:21]
  wire  _T_75; // @[LZD.scala 39:30]
  wire  _T_76; // @[LZD.scala 39:27]
  wire  _T_77; // @[LZD.scala 39:25]
  wire [1:0] _T_78; // @[Cat.scala 29:58]
  wire  _T_79; // @[Shift.scala 12:21]
  wire  _T_80; // @[Shift.scala 12:21]
  wire  _T_81; // @[LZD.scala 49:16]
  wire  _T_82; // @[LZD.scala 49:27]
  wire  _T_83; // @[LZD.scala 49:25]
  wire  _T_84; // @[LZD.scala 49:47]
  wire  _T_85; // @[LZD.scala 49:59]
  wire  _T_86; // @[LZD.scala 49:35]
  wire [2:0] _T_88; // @[Cat.scala 29:58]
  wire  _T_89; // @[LZD.scala 44:32]
  wire  _T_91; // @[Shift.scala 12:21]
  wire [1:0] _T_93; // @[Cat.scala 29:58]
  wire [1:0] _T_94; // @[LZD.scala 55:32]
  wire [1:0] _T_95; // @[LZD.scala 55:20]
  wire [2:0] _T_96; // @[Cat.scala 29:58]
  wire  _T_97; // @[Shift.scala 12:21]
  wire [2:0] _T_99; // @[LZD.scala 55:32]
  wire [2:0] _T_100; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [3:0] shiftValue; // @[FMAEnc.scala 37:24]
  wire [11:0] _T_101; // @[FMAEnc.scala 38:41]
  wire  _T_102; // @[Shift.scala 16:24]
  wire  _T_104; // @[Shift.scala 12:21]
  wire [3:0] _T_105; // @[Shift.scala 64:52]
  wire [11:0] _T_107; // @[Cat.scala 29:58]
  wire [11:0] _T_108; // @[Shift.scala 64:27]
  wire [2:0] _T_109; // @[Shift.scala 66:70]
  wire  _T_110; // @[Shift.scala 12:21]
  wire [7:0] _T_111; // @[Shift.scala 64:52]
  wire [11:0] _T_113; // @[Cat.scala 29:58]
  wire [11:0] _T_114; // @[Shift.scala 64:27]
  wire [1:0] _T_115; // @[Shift.scala 66:70]
  wire  _T_116; // @[Shift.scala 12:21]
  wire [9:0] _T_117; // @[Shift.scala 64:52]
  wire [11:0] _T_119; // @[Cat.scala 29:58]
  wire [11:0] _T_120; // @[Shift.scala 64:27]
  wire  _T_121; // @[Shift.scala 66:70]
  wire [10:0] _T_123; // @[Shift.scala 64:52]
  wire [11:0] _T_124; // @[Cat.scala 29:58]
  wire [11:0] _T_125; // @[Shift.scala 64:27]
  wire [11:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [3:0] _T_127; // @[FMAEnc.scala 41:39]
  wire [3:0] _T_128; // @[FMAEnc.scala 41:39]
  wire [4:0] _T_129; // @[Cat.scala 29:58]
  wire [4:0] _T_130; // @[FMAEnc.scala 41:64]
  wire [4:0] _GEN_2; // @[FMAEnc.scala 41:45]
  wire [4:0] _T_132; // @[FMAEnc.scala 41:45]
  wire [4:0] sumScale; // @[FMAEnc.scala 41:45]
  wire [4:0] sumFrac; // @[FMAEnc.scala 42:41]
  wire [6:0] grsTmp; // @[FMAEnc.scala 45:41]
  wire [1:0] _T_133; // @[FMAEnc.scala 48:40]
  wire [4:0] _T_134; // @[FMAEnc.scala 48:56]
  wire  _T_135; // @[FMAEnc.scala 48:60]
  wire  underflow; // @[FMAEnc.scala 55:32]
  wire  overflow; // @[FMAEnc.scala 56:32]
  wire  _T_136; // @[FMAEnc.scala 65:35]
  wire  decF_isZero; // @[FMAEnc.scala 65:20]
  wire [4:0] _T_138; // @[Mux.scala 87:16]
  wire [4:0] _T_139; // @[Mux.scala 87:16]
  wire [3:0] _GEN_3; // @[FMAEnc.scala 62:18 FMAEnc.scala 68:17]
  wire [3:0] decF_scale; // @[FMAEnc.scala 62:18 FMAEnc.scala 68:17]
  wire  _T_141; // @[convert.scala 49:36]
  wire [3:0] _T_143; // @[convert.scala 50:36]
  wire [3:0] _T_144; // @[convert.scala 50:36]
  wire [3:0] _T_145; // @[convert.scala 50:28]
  wire  _T_146; // @[convert.scala 51:31]
  wire  _T_147; // @[convert.scala 53:34]
  wire [9:0] _T_150; // @[Cat.scala 29:58]
  wire [3:0] _T_151; // @[Shift.scala 39:17]
  wire  _T_152; // @[Shift.scala 39:24]
  wire [1:0] _T_154; // @[Shift.scala 90:30]
  wire [7:0] _T_155; // @[Shift.scala 90:48]
  wire  _T_156; // @[Shift.scala 90:57]
  wire [1:0] _GEN_4; // @[Shift.scala 90:39]
  wire [1:0] _T_157; // @[Shift.scala 90:39]
  wire  _T_158; // @[Shift.scala 12:21]
  wire  _T_159; // @[Shift.scala 12:21]
  wire [7:0] _T_161; // @[Bitwise.scala 71:12]
  wire [9:0] _T_162; // @[Cat.scala 29:58]
  wire [9:0] _T_163; // @[Shift.scala 91:22]
  wire [2:0] _T_164; // @[Shift.scala 92:77]
  wire [5:0] _T_165; // @[Shift.scala 90:30]
  wire [3:0] _T_166; // @[Shift.scala 90:48]
  wire  _T_167; // @[Shift.scala 90:57]
  wire [5:0] _GEN_5; // @[Shift.scala 90:39]
  wire [5:0] _T_168; // @[Shift.scala 90:39]
  wire  _T_169; // @[Shift.scala 12:21]
  wire  _T_170; // @[Shift.scala 12:21]
  wire [3:0] _T_172; // @[Bitwise.scala 71:12]
  wire [9:0] _T_173; // @[Cat.scala 29:58]
  wire [9:0] _T_174; // @[Shift.scala 91:22]
  wire [1:0] _T_175; // @[Shift.scala 92:77]
  wire [7:0] _T_176; // @[Shift.scala 90:30]
  wire [1:0] _T_177; // @[Shift.scala 90:48]
  wire  _T_178; // @[Shift.scala 90:57]
  wire [7:0] _GEN_6; // @[Shift.scala 90:39]
  wire [7:0] _T_179; // @[Shift.scala 90:39]
  wire  _T_180; // @[Shift.scala 12:21]
  wire  _T_181; // @[Shift.scala 12:21]
  wire [1:0] _T_183; // @[Bitwise.scala 71:12]
  wire [9:0] _T_184; // @[Cat.scala 29:58]
  wire [9:0] _T_185; // @[Shift.scala 91:22]
  wire  _T_186; // @[Shift.scala 92:77]
  wire [8:0] _T_187; // @[Shift.scala 90:30]
  wire  _T_188; // @[Shift.scala 90:48]
  wire [8:0] _GEN_7; // @[Shift.scala 90:39]
  wire [8:0] _T_190; // @[Shift.scala 90:39]
  wire  _T_192; // @[Shift.scala 12:21]
  wire [9:0] _T_193; // @[Cat.scala 29:58]
  wire [9:0] _T_194; // @[Shift.scala 91:22]
  wire [9:0] _T_197; // @[Bitwise.scala 71:12]
  wire [9:0] _T_198; // @[Shift.scala 39:10]
  wire  _T_199; // @[convert.scala 55:31]
  wire  _T_200; // @[convert.scala 56:31]
  wire  _T_201; // @[convert.scala 57:31]
  wire  _T_202; // @[convert.scala 58:31]
  wire [6:0] _T_203; // @[convert.scala 59:69]
  wire  _T_204; // @[convert.scala 59:81]
  wire  _T_205; // @[convert.scala 59:50]
  wire  _T_207; // @[convert.scala 60:81]
  wire  _T_208; // @[convert.scala 61:44]
  wire  _T_209; // @[convert.scala 61:52]
  wire  _T_210; // @[convert.scala 61:36]
  wire  _T_211; // @[convert.scala 62:63]
  wire  _T_212; // @[convert.scala 62:103]
  wire  _T_213; // @[convert.scala 62:60]
  wire [6:0] _GEN_8; // @[convert.scala 63:56]
  wire [6:0] _T_216; // @[convert.scala 63:56]
  wire [7:0] _T_217; // @[Cat.scala 29:58]
  reg  _T_221; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [7:0] _T_225; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  assign _T = io_signSumSig[13:1]; // @[FMAEnc.scala 35:36]
  assign _T_1 = io_signSumSig[12:0]; // @[FMAEnc.scala 35:74]
  assign sumXor = _T ^ _T_1; // @[FMAEnc.scala 35:54]
  assign _T_2 = sumXor[12:5]; // @[LZD.scala 43:32]
  assign _T_3 = _T_2[7:4]; // @[LZD.scala 43:32]
  assign _T_4 = _T_3[3:2]; // @[LZD.scala 43:32]
  assign _T_5 = _T_4 != 2'h0; // @[LZD.scala 39:14]
  assign _T_6 = _T_4[1]; // @[LZD.scala 39:21]
  assign _T_7 = _T_4[0]; // @[LZD.scala 39:30]
  assign _T_8 = ~ _T_7; // @[LZD.scala 39:27]
  assign _T_9 = _T_6 | _T_8; // @[LZD.scala 39:25]
  assign _T_10 = {_T_5,_T_9}; // @[Cat.scala 29:58]
  assign _T_11 = _T_3[1:0]; // @[LZD.scala 44:32]
  assign _T_12 = _T_11 != 2'h0; // @[LZD.scala 39:14]
  assign _T_13 = _T_11[1]; // @[LZD.scala 39:21]
  assign _T_14 = _T_11[0]; // @[LZD.scala 39:30]
  assign _T_15 = ~ _T_14; // @[LZD.scala 39:27]
  assign _T_16 = _T_13 | _T_15; // @[LZD.scala 39:25]
  assign _T_17 = {_T_12,_T_16}; // @[Cat.scala 29:58]
  assign _T_18 = _T_10[1]; // @[Shift.scala 12:21]
  assign _T_19 = _T_17[1]; // @[Shift.scala 12:21]
  assign _T_20 = _T_18 | _T_19; // @[LZD.scala 49:16]
  assign _T_21 = ~ _T_19; // @[LZD.scala 49:27]
  assign _T_22 = _T_18 | _T_21; // @[LZD.scala 49:25]
  assign _T_23 = _T_10[0:0]; // @[LZD.scala 49:47]
  assign _T_24 = _T_17[0:0]; // @[LZD.scala 49:59]
  assign _T_25 = _T_18 ? _T_23 : _T_24; // @[LZD.scala 49:35]
  assign _T_27 = {_T_20,_T_22,_T_25}; // @[Cat.scala 29:58]
  assign _T_28 = _T_2[3:0]; // @[LZD.scala 44:32]
  assign _T_29 = _T_28[3:2]; // @[LZD.scala 43:32]
  assign _T_30 = _T_29 != 2'h0; // @[LZD.scala 39:14]
  assign _T_31 = _T_29[1]; // @[LZD.scala 39:21]
  assign _T_32 = _T_29[0]; // @[LZD.scala 39:30]
  assign _T_33 = ~ _T_32; // @[LZD.scala 39:27]
  assign _T_34 = _T_31 | _T_33; // @[LZD.scala 39:25]
  assign _T_35 = {_T_30,_T_34}; // @[Cat.scala 29:58]
  assign _T_36 = _T_28[1:0]; // @[LZD.scala 44:32]
  assign _T_37 = _T_36 != 2'h0; // @[LZD.scala 39:14]
  assign _T_38 = _T_36[1]; // @[LZD.scala 39:21]
  assign _T_39 = _T_36[0]; // @[LZD.scala 39:30]
  assign _T_40 = ~ _T_39; // @[LZD.scala 39:27]
  assign _T_41 = _T_38 | _T_40; // @[LZD.scala 39:25]
  assign _T_42 = {_T_37,_T_41}; // @[Cat.scala 29:58]
  assign _T_43 = _T_35[1]; // @[Shift.scala 12:21]
  assign _T_44 = _T_42[1]; // @[Shift.scala 12:21]
  assign _T_45 = _T_43 | _T_44; // @[LZD.scala 49:16]
  assign _T_46 = ~ _T_44; // @[LZD.scala 49:27]
  assign _T_47 = _T_43 | _T_46; // @[LZD.scala 49:25]
  assign _T_48 = _T_35[0:0]; // @[LZD.scala 49:47]
  assign _T_49 = _T_42[0:0]; // @[LZD.scala 49:59]
  assign _T_50 = _T_43 ? _T_48 : _T_49; // @[LZD.scala 49:35]
  assign _T_52 = {_T_45,_T_47,_T_50}; // @[Cat.scala 29:58]
  assign _T_53 = _T_27[2]; // @[Shift.scala 12:21]
  assign _T_54 = _T_52[2]; // @[Shift.scala 12:21]
  assign _T_55 = _T_53 | _T_54; // @[LZD.scala 49:16]
  assign _T_56 = ~ _T_54; // @[LZD.scala 49:27]
  assign _T_57 = _T_53 | _T_56; // @[LZD.scala 49:25]
  assign _T_58 = _T_27[1:0]; // @[LZD.scala 49:47]
  assign _T_59 = _T_52[1:0]; // @[LZD.scala 49:59]
  assign _T_60 = _T_53 ? _T_58 : _T_59; // @[LZD.scala 49:35]
  assign _T_62 = {_T_55,_T_57,_T_60}; // @[Cat.scala 29:58]
  assign _T_63 = sumXor[4:0]; // @[LZD.scala 44:32]
  assign _T_64 = _T_63[4:1]; // @[LZD.scala 43:32]
  assign _T_65 = _T_64[3:2]; // @[LZD.scala 43:32]
  assign _T_66 = _T_65 != 2'h0; // @[LZD.scala 39:14]
  assign _T_67 = _T_65[1]; // @[LZD.scala 39:21]
  assign _T_68 = _T_65[0]; // @[LZD.scala 39:30]
  assign _T_69 = ~ _T_68; // @[LZD.scala 39:27]
  assign _T_70 = _T_67 | _T_69; // @[LZD.scala 39:25]
  assign _T_71 = {_T_66,_T_70}; // @[Cat.scala 29:58]
  assign _T_72 = _T_64[1:0]; // @[LZD.scala 44:32]
  assign _T_73 = _T_72 != 2'h0; // @[LZD.scala 39:14]
  assign _T_74 = _T_72[1]; // @[LZD.scala 39:21]
  assign _T_75 = _T_72[0]; // @[LZD.scala 39:30]
  assign _T_76 = ~ _T_75; // @[LZD.scala 39:27]
  assign _T_77 = _T_74 | _T_76; // @[LZD.scala 39:25]
  assign _T_78 = {_T_73,_T_77}; // @[Cat.scala 29:58]
  assign _T_79 = _T_71[1]; // @[Shift.scala 12:21]
  assign _T_80 = _T_78[1]; // @[Shift.scala 12:21]
  assign _T_81 = _T_79 | _T_80; // @[LZD.scala 49:16]
  assign _T_82 = ~ _T_80; // @[LZD.scala 49:27]
  assign _T_83 = _T_79 | _T_82; // @[LZD.scala 49:25]
  assign _T_84 = _T_71[0:0]; // @[LZD.scala 49:47]
  assign _T_85 = _T_78[0:0]; // @[LZD.scala 49:59]
  assign _T_86 = _T_79 ? _T_84 : _T_85; // @[LZD.scala 49:35]
  assign _T_88 = {_T_81,_T_83,_T_86}; // @[Cat.scala 29:58]
  assign _T_89 = _T_63[0:0]; // @[LZD.scala 44:32]
  assign _T_91 = _T_88[2]; // @[Shift.scala 12:21]
  assign _T_93 = {1'h1,_T_89}; // @[Cat.scala 29:58]
  assign _T_94 = _T_88[1:0]; // @[LZD.scala 55:32]
  assign _T_95 = _T_91 ? _T_94 : _T_93; // @[LZD.scala 55:20]
  assign _T_96 = {_T_91,_T_95}; // @[Cat.scala 29:58]
  assign _T_97 = _T_62[3]; // @[Shift.scala 12:21]
  assign _T_99 = _T_62[2:0]; // @[LZD.scala 55:32]
  assign _T_100 = _T_97 ? _T_99 : _T_96; // @[LZD.scala 55:20]
  assign sumLZD = {_T_97,_T_100}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[FMAEnc.scala 37:24]
  assign _T_101 = io_signSumSig[11:0]; // @[FMAEnc.scala 38:41]
  assign _T_102 = shiftValue < 4'hc; // @[Shift.scala 16:24]
  assign _T_104 = shiftValue[3]; // @[Shift.scala 12:21]
  assign _T_105 = _T_101[3:0]; // @[Shift.scala 64:52]
  assign _T_107 = {_T_105,8'h0}; // @[Cat.scala 29:58]
  assign _T_108 = _T_104 ? _T_107 : _T_101; // @[Shift.scala 64:27]
  assign _T_109 = shiftValue[2:0]; // @[Shift.scala 66:70]
  assign _T_110 = _T_109[2]; // @[Shift.scala 12:21]
  assign _T_111 = _T_108[7:0]; // @[Shift.scala 64:52]
  assign _T_113 = {_T_111,4'h0}; // @[Cat.scala 29:58]
  assign _T_114 = _T_110 ? _T_113 : _T_108; // @[Shift.scala 64:27]
  assign _T_115 = _T_109[1:0]; // @[Shift.scala 66:70]
  assign _T_116 = _T_115[1]; // @[Shift.scala 12:21]
  assign _T_117 = _T_114[9:0]; // @[Shift.scala 64:52]
  assign _T_119 = {_T_117,2'h0}; // @[Cat.scala 29:58]
  assign _T_120 = _T_116 ? _T_119 : _T_114; // @[Shift.scala 64:27]
  assign _T_121 = _T_115[0:0]; // @[Shift.scala 66:70]
  assign _T_123 = _T_120[10:0]; // @[Shift.scala 64:52]
  assign _T_124 = {_T_123,1'h0}; // @[Cat.scala 29:58]
  assign _T_125 = _T_121 ? _T_124 : _T_120; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_102 ? _T_125 : 12'h0; // @[Shift.scala 16:10]
  assign _T_127 = $signed(io_greaterScale) + $signed(4'sh2); // @[FMAEnc.scala 41:39]
  assign _T_128 = $signed(_T_127); // @[FMAEnc.scala 41:39]
  assign _T_129 = {1'h1,_T_97,_T_100}; // @[Cat.scala 29:58]
  assign _T_130 = $signed(_T_129); // @[FMAEnc.scala 41:64]
  assign _GEN_2 = {{1{_T_128[3]}},_T_128}; // @[FMAEnc.scala 41:45]
  assign _T_132 = $signed(_GEN_2) + $signed(_T_130); // @[FMAEnc.scala 41:45]
  assign sumScale = $signed(_T_132); // @[FMAEnc.scala 41:45]
  assign sumFrac = normalFracTmp[11:7]; // @[FMAEnc.scala 42:41]
  assign grsTmp = normalFracTmp[6:0]; // @[FMAEnc.scala 45:41]
  assign _T_133 = grsTmp[6:5]; // @[FMAEnc.scala 48:40]
  assign _T_134 = grsTmp[4:0]; // @[FMAEnc.scala 48:56]
  assign _T_135 = _T_134 != 5'h0; // @[FMAEnc.scala 48:60]
  assign underflow = $signed(sumScale) < $signed(-5'sh7); // @[FMAEnc.scala 55:32]
  assign overflow = $signed(sumScale) > $signed(5'sh6); // @[FMAEnc.scala 56:32]
  assign _T_136 = io_signSumSig != 14'h0; // @[FMAEnc.scala 65:35]
  assign decF_isZero = ~ _T_136; // @[FMAEnc.scala 65:20]
  assign _T_138 = underflow ? $signed(-5'sh7) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_139 = overflow ? $signed(5'sh6) : $signed(_T_138); // @[Mux.scala 87:16]
  assign _GEN_3 = _T_139[3:0]; // @[FMAEnc.scala 62:18 FMAEnc.scala 68:17]
  assign decF_scale = $signed(_GEN_3); // @[FMAEnc.scala 62:18 FMAEnc.scala 68:17]
  assign _T_141 = decF_scale[3:3]; // @[convert.scala 49:36]
  assign _T_143 = ~ decF_scale; // @[convert.scala 50:36]
  assign _T_144 = $signed(_T_143); // @[convert.scala 50:36]
  assign _T_145 = _T_141 ? $signed(_T_144) : $signed(decF_scale); // @[convert.scala 50:28]
  assign _T_146 = _T_141 ^ io_sumSign; // @[convert.scala 51:31]
  assign _T_147 = ~ _T_146; // @[convert.scala 53:34]
  assign _T_150 = {_T_147,_T_146,sumFrac,_T_133,_T_135}; // @[Cat.scala 29:58]
  assign _T_151 = $unsigned(_T_145); // @[Shift.scala 39:17]
  assign _T_152 = _T_151 < 4'ha; // @[Shift.scala 39:24]
  assign _T_154 = _T_150[9:8]; // @[Shift.scala 90:30]
  assign _T_155 = _T_150[7:0]; // @[Shift.scala 90:48]
  assign _T_156 = _T_155 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_4 = {{1'd0}, _T_156}; // @[Shift.scala 90:39]
  assign _T_157 = _T_154 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_158 = _T_151[3]; // @[Shift.scala 12:21]
  assign _T_159 = _T_150[9]; // @[Shift.scala 12:21]
  assign _T_161 = _T_159 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_162 = {_T_161,_T_157}; // @[Cat.scala 29:58]
  assign _T_163 = _T_158 ? _T_162 : _T_150; // @[Shift.scala 91:22]
  assign _T_164 = _T_151[2:0]; // @[Shift.scala 92:77]
  assign _T_165 = _T_163[9:4]; // @[Shift.scala 90:30]
  assign _T_166 = _T_163[3:0]; // @[Shift.scala 90:48]
  assign _T_167 = _T_166 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{5'd0}, _T_167}; // @[Shift.scala 90:39]
  assign _T_168 = _T_165 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_169 = _T_164[2]; // @[Shift.scala 12:21]
  assign _T_170 = _T_163[9]; // @[Shift.scala 12:21]
  assign _T_172 = _T_170 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_173 = {_T_172,_T_168}; // @[Cat.scala 29:58]
  assign _T_174 = _T_169 ? _T_173 : _T_163; // @[Shift.scala 91:22]
  assign _T_175 = _T_164[1:0]; // @[Shift.scala 92:77]
  assign _T_176 = _T_174[9:2]; // @[Shift.scala 90:30]
  assign _T_177 = _T_174[1:0]; // @[Shift.scala 90:48]
  assign _T_178 = _T_177 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{7'd0}, _T_178}; // @[Shift.scala 90:39]
  assign _T_179 = _T_176 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_180 = _T_175[1]; // @[Shift.scala 12:21]
  assign _T_181 = _T_174[9]; // @[Shift.scala 12:21]
  assign _T_183 = _T_181 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_184 = {_T_183,_T_179}; // @[Cat.scala 29:58]
  assign _T_185 = _T_180 ? _T_184 : _T_174; // @[Shift.scala 91:22]
  assign _T_186 = _T_175[0:0]; // @[Shift.scala 92:77]
  assign _T_187 = _T_185[9:1]; // @[Shift.scala 90:30]
  assign _T_188 = _T_185[0:0]; // @[Shift.scala 90:48]
  assign _GEN_7 = {{8'd0}, _T_188}; // @[Shift.scala 90:39]
  assign _T_190 = _T_187 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_192 = _T_185[9]; // @[Shift.scala 12:21]
  assign _T_193 = {_T_192,_T_190}; // @[Cat.scala 29:58]
  assign _T_194 = _T_186 ? _T_193 : _T_185; // @[Shift.scala 91:22]
  assign _T_197 = _T_159 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_198 = _T_152 ? _T_194 : _T_197; // @[Shift.scala 39:10]
  assign _T_199 = _T_198[3]; // @[convert.scala 55:31]
  assign _T_200 = _T_198[2]; // @[convert.scala 56:31]
  assign _T_201 = _T_198[1]; // @[convert.scala 57:31]
  assign _T_202 = _T_198[0]; // @[convert.scala 58:31]
  assign _T_203 = _T_198[9:3]; // @[convert.scala 59:69]
  assign _T_204 = _T_203 != 7'h0; // @[convert.scala 59:81]
  assign _T_205 = ~ _T_204; // @[convert.scala 59:50]
  assign _T_207 = _T_203 == 7'h7f; // @[convert.scala 60:81]
  assign _T_208 = _T_199 | _T_201; // @[convert.scala 61:44]
  assign _T_209 = _T_208 | _T_202; // @[convert.scala 61:52]
  assign _T_210 = _T_200 & _T_209; // @[convert.scala 61:36]
  assign _T_211 = ~ _T_207; // @[convert.scala 62:63]
  assign _T_212 = _T_211 & _T_210; // @[convert.scala 62:103]
  assign _T_213 = _T_205 | _T_212; // @[convert.scala 62:60]
  assign _GEN_8 = {{6'd0}, _T_213}; // @[convert.scala 63:56]
  assign _T_216 = _T_203 + _GEN_8; // @[convert.scala 63:56]
  assign _T_217 = {io_sumSign,_T_216}; // @[Cat.scala 29:58]
  assign io_F = _T_225; // @[FMAEnc.scala 85:15]
  assign io_outValid = _T_221; // @[FMAEnc.scala 84:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_221 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_225 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_221 <= 1'h0;
    end else begin
      _T_221 <= io_inValid_phase2;
    end
    if (io_inValid_phase2) begin
      if (io_outIsNaR_phase2) begin
        _T_225 <= 8'h80;
      end else begin
        if (decF_isZero) begin
          _T_225 <= 8'h0;
        end else begin
          _T_225 <= _T_217;
        end
      end
    end
  end
endmodule
