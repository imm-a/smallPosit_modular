module PositDivSqrter7_0(
  input        clock,
  input        reset,
  output       io_inReady,
  input        io_inValid,
  input        io_sqrtOp,
  input  [6:0] io_A,
  input  [6:0] io_B,
  output       io_diviValid,
  output       io_sqrtValid,
  output       io_invalidExc,
  output [6:0] io_Q
);
  reg [3:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [4:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg [3:0] fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [10:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [10:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [4:0] _T_4; // @[convert.scala 19:24]
  wire [4:0] _T_5; // @[convert.scala 19:43]
  wire [4:0] _T_6; // @[convert.scala 19:39]
  wire [3:0] _T_7; // @[LZD.scala 43:32]
  wire [1:0] _T_8; // @[LZD.scala 43:32]
  wire  _T_9; // @[LZD.scala 39:14]
  wire  _T_10; // @[LZD.scala 39:21]
  wire  _T_11; // @[LZD.scala 39:30]
  wire  _T_12; // @[LZD.scala 39:27]
  wire  _T_13; // @[LZD.scala 39:25]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [1:0] _T_15; // @[LZD.scala 44:32]
  wire  _T_16; // @[LZD.scala 39:14]
  wire  _T_17; // @[LZD.scala 39:21]
  wire  _T_18; // @[LZD.scala 39:30]
  wire  _T_19; // @[LZD.scala 39:27]
  wire  _T_20; // @[LZD.scala 39:25]
  wire [1:0] _T_21; // @[Cat.scala 29:58]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[LZD.scala 49:16]
  wire  _T_25; // @[LZD.scala 49:27]
  wire  _T_26; // @[LZD.scala 49:25]
  wire  _T_27; // @[LZD.scala 49:47]
  wire  _T_28; // @[LZD.scala 49:59]
  wire  _T_29; // @[LZD.scala 49:35]
  wire [2:0] _T_31; // @[Cat.scala 29:58]
  wire  _T_32; // @[LZD.scala 44:32]
  wire  _T_34; // @[Shift.scala 12:21]
  wire [1:0] _T_36; // @[Cat.scala 29:58]
  wire [1:0] _T_37; // @[LZD.scala 55:32]
  wire [1:0] _T_38; // @[LZD.scala 55:20]
  wire [2:0] _T_39; // @[Cat.scala 29:58]
  wire [2:0] _T_40; // @[convert.scala 21:22]
  wire [3:0] _T_41; // @[convert.scala 22:36]
  wire  _T_42; // @[Shift.scala 16:24]
  wire [1:0] _T_43; // @[Shift.scala 17:37]
  wire  _T_44; // @[Shift.scala 12:21]
  wire [1:0] _T_45; // @[Shift.scala 64:52]
  wire [3:0] _T_47; // @[Cat.scala 29:58]
  wire [3:0] _T_48; // @[Shift.scala 64:27]
  wire  _T_49; // @[Shift.scala 66:70]
  wire [2:0] _T_51; // @[Shift.scala 64:52]
  wire [3:0] _T_52; // @[Cat.scala 29:58]
  wire [3:0] _T_53; // @[Shift.scala 64:27]
  wire [3:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_57; // @[convert.scala 25:26]
  wire [2:0] _T_59; // @[convert.scala 25:42]
  wire [3:0] _T_60; // @[Cat.scala 29:58]
  wire [5:0] _T_62; // @[convert.scala 29:56]
  wire  _T_63; // @[convert.scala 29:60]
  wire  _T_64; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_67; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [3:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_76; // @[convert.scala 18:24]
  wire  _T_77; // @[convert.scala 18:40]
  wire  _T_78; // @[convert.scala 18:36]
  wire [4:0] _T_79; // @[convert.scala 19:24]
  wire [4:0] _T_80; // @[convert.scala 19:43]
  wire [4:0] _T_81; // @[convert.scala 19:39]
  wire [3:0] _T_82; // @[LZD.scala 43:32]
  wire [1:0] _T_83; // @[LZD.scala 43:32]
  wire  _T_84; // @[LZD.scala 39:14]
  wire  _T_85; // @[LZD.scala 39:21]
  wire  _T_86; // @[LZD.scala 39:30]
  wire  _T_87; // @[LZD.scala 39:27]
  wire  _T_88; // @[LZD.scala 39:25]
  wire [1:0] _T_89; // @[Cat.scala 29:58]
  wire [1:0] _T_90; // @[LZD.scala 44:32]
  wire  _T_91; // @[LZD.scala 39:14]
  wire  _T_92; // @[LZD.scala 39:21]
  wire  _T_93; // @[LZD.scala 39:30]
  wire  _T_94; // @[LZD.scala 39:27]
  wire  _T_95; // @[LZD.scala 39:25]
  wire [1:0] _T_96; // @[Cat.scala 29:58]
  wire  _T_97; // @[Shift.scala 12:21]
  wire  _T_98; // @[Shift.scala 12:21]
  wire  _T_99; // @[LZD.scala 49:16]
  wire  _T_100; // @[LZD.scala 49:27]
  wire  _T_101; // @[LZD.scala 49:25]
  wire  _T_102; // @[LZD.scala 49:47]
  wire  _T_103; // @[LZD.scala 49:59]
  wire  _T_104; // @[LZD.scala 49:35]
  wire [2:0] _T_106; // @[Cat.scala 29:58]
  wire  _T_107; // @[LZD.scala 44:32]
  wire  _T_109; // @[Shift.scala 12:21]
  wire [1:0] _T_111; // @[Cat.scala 29:58]
  wire [1:0] _T_112; // @[LZD.scala 55:32]
  wire [1:0] _T_113; // @[LZD.scala 55:20]
  wire [2:0] _T_114; // @[Cat.scala 29:58]
  wire [2:0] _T_115; // @[convert.scala 21:22]
  wire [3:0] _T_116; // @[convert.scala 22:36]
  wire  _T_117; // @[Shift.scala 16:24]
  wire [1:0] _T_118; // @[Shift.scala 17:37]
  wire  _T_119; // @[Shift.scala 12:21]
  wire [1:0] _T_120; // @[Shift.scala 64:52]
  wire [3:0] _T_122; // @[Cat.scala 29:58]
  wire [3:0] _T_123; // @[Shift.scala 64:27]
  wire  _T_124; // @[Shift.scala 66:70]
  wire [2:0] _T_126; // @[Shift.scala 64:52]
  wire [3:0] _T_127; // @[Cat.scala 29:58]
  wire [3:0] _T_128; // @[Shift.scala 64:27]
  wire [3:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_132; // @[convert.scala 25:26]
  wire [2:0] _T_134; // @[convert.scala 25:42]
  wire [3:0] _T_135; // @[Cat.scala 29:58]
  wire [5:0] _T_137; // @[convert.scala 29:56]
  wire  _T_138; // @[convert.scala 29:60]
  wire  _T_139; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_142; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [3:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_151; // @[Bitwise.scala 71:12]
  wire  _T_152; // @[PositDivisionSqrt.scala 80:40]
  wire [10:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_155; // @[PositDivisionSqrt.scala 82:31]
  wire [10:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_158; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_159; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_160; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_161; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_162; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_163; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_164; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_165; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_166; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_167; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [4:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_170; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_171; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_172; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_173; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_174; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_175; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_176; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_177; // @[PositDivisionSqrt.scala 117:30]
  wire [3:0] _T_179; // @[PositDivisionSqrt.scala 119:26]
  wire [3:0] _T_180; // @[PositDivisionSqrt.scala 118:20]
  wire [3:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [3:0] _T_181; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_183; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_184; // @[PositDivisionSqrt.scala 123:27]
  wire [3:0] _T_186; // @[PositDivisionSqrt.scala 123:52]
  wire [3:0] _T_187; // @[PositDivisionSqrt.scala 123:20]
  wire [3:0] _T_188; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_190; // @[PositDivisionSqrt.scala 124:27]
  wire [3:0] _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _T_192; // @[PositDivisionSqrt.scala 123:64]
  wire [2:0] _T_193; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_195; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_196; // @[PositDivisionSqrt.scala 137:28]
  wire [15:0] _T_197; // @[PositDivisionSqrt.scala 146:22]
  wire [13:0] _T_198; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_199; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_200; // @[PositDivisionSqrt.scala 148:23]
  wire [10:0] _T_201; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_202; // @[PositDivisionSqrt.scala 149:23]
  wire [11:0] _T_203; // @[PositDivisionSqrt.scala 149:46]
  wire [10:0] _T_204; // @[PositDivisionSqrt.scala 149:56]
  wire [10:0] _T_205; // @[PositDivisionSqrt.scala 149:16]
  wire [10:0] _T_206; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_207; // @[PositDivisionSqrt.scala 150:17]
  wire [10:0] _T_208; // @[PositDivisionSqrt.scala 150:16]
  wire [10:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_210; // @[PositDivisionSqrt.scala 152:29]
  wire [10:0] _T_211; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_212; // @[PositDivisionSqrt.scala 153:29]
  wire [7:0] _T_213; // @[PositDivisionSqrt.scala 153:22]
  wire [10:0] _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  wire [10:0] _T_214; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_216; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_217; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_218; // @[PositDivisionSqrt.scala 154:57]
  wire [10:0] _T_221; // @[Cat.scala 29:58]
  wire [10:0] _T_222; // @[PositDivisionSqrt.scala 154:22]
  wire [10:0] _T_223; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_225; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_226; // @[PositDivisionSqrt.scala 156:83]
  wire [6:0] _T_228; // @[Bitwise.scala 71:12]
  wire [9:0] bitMask; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  wire [9:0] _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  wire [9:0] _T_229; // @[PositDivisionSqrt.scala 156:53]
  wire [10:0] _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  wire [10:0] _T_230; // @[PositDivisionSqrt.scala 155:51]
  wire [8:0] _T_231; // @[PositDivisionSqrt.scala 157:53]
  wire [10:0] _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  wire [10:0] _T_232; // @[PositDivisionSqrt.scala 156:89]
  wire [10:0] _T_233; // @[PositDivisionSqrt.scala 155:22]
  wire [10:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_235; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_236; // @[PositDivisionSqrt.scala 162:40]
  wire [10:0] _T_239; // @[PositDivisionSqrt.scala 163:97]
  wire [10:0] _T_241; // @[PositDivisionSqrt.scala 164:97]
  wire [10:0] _T_242; // @[PositDivisionSqrt.scala 161:92]
  wire [11:0] _T_247; // @[PositDivisionSqrt.scala 168:98]
  wire [10:0] _T_248; // @[PositDivisionSqrt.scala 168:108]
  wire [10:0] _T_250; // @[PositDivisionSqrt.scala 168:112]
  wire [10:0] _T_254; // @[PositDivisionSqrt.scala 169:112]
  wire [10:0] _T_255; // @[PositDivisionSqrt.scala 166:26]
  wire [10:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_256; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_257; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_259; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_260; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_261; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_262; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_263; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_265; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_266; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_267; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_268; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_269; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_272; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_273; // @[PositDivisionSqrt.scala 187:28]
  wire [10:0] _T_276; // @[PositDivisionSqrt.scala 188:47]
  wire [10:0] _T_277; // @[PositDivisionSqrt.scala 188:18]
  wire [8:0] _T_279; // @[PositDivisionSqrt.scala 189:18]
  wire [10:0] _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  wire [10:0] _T_280; // @[PositDivisionSqrt.scala 188:78]
  wire [10:0] _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  wire [10:0] _T_282; // @[PositDivisionSqrt.scala 190:47]
  wire [10:0] _T_283; // @[PositDivisionSqrt.scala 190:18]
  wire [10:0] _T_284; // @[PositDivisionSqrt.scala 189:78]
  wire [1:0] _T_286; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [10:0] _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  wire [10:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire [3:0] _T_289; // @[PositDivisionSqrt.scala 200:97]
  wire [3:0] _T_290; // @[PositDivisionSqrt.scala 201:97]
  wire [3:0] realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_291; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_292; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_293; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  _T_295; // @[PositDivisionSqrt.scala 206:56]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_296; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_297; // @[Cat.scala 29:58]
  wire [2:0] _T_298; // @[PositDivisionSqrt.scala 209:63]
  wire [4:0] _GEN_18; // @[PositDivisionSqrt.scala 209:31]
  wire [4:0] _T_300; // @[PositDivisionSqrt.scala 209:31]
  wire [4:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [4:0] _T_302; // @[Mux.scala 87:16]
  wire [4:0] _T_303; // @[Mux.scala 87:16]
  wire [2:0] _T_304; // @[PositDivisionSqrt.scala 224:48]
  wire [2:0] _T_305; // @[PositDivisionSqrt.scala 224:64]
  wire [2:0] decQ_grs; // @[PositDivisionSqrt.scala 224:23]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [3:0] _GEN_19; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [3:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire  _T_312; // @[convert.scala 49:36]
  wire [3:0] _T_314; // @[convert.scala 50:36]
  wire [3:0] _T_315; // @[convert.scala 50:36]
  wire [3:0] _T_316; // @[convert.scala 50:28]
  wire  _T_317; // @[convert.scala 51:31]
  wire  _T_318; // @[convert.scala 53:34]
  wire [8:0] _T_321; // @[Cat.scala 29:58]
  wire [3:0] _T_322; // @[Shift.scala 39:17]
  wire  _T_323; // @[Shift.scala 39:24]
  wire  _T_325; // @[Shift.scala 90:30]
  wire [7:0] _T_326; // @[Shift.scala 90:48]
  wire  _T_327; // @[Shift.scala 90:57]
  wire  _T_328; // @[Shift.scala 90:39]
  wire  _T_329; // @[Shift.scala 12:21]
  wire  _T_330; // @[Shift.scala 12:21]
  wire [7:0] _T_332; // @[Bitwise.scala 71:12]
  wire [8:0] _T_333; // @[Cat.scala 29:58]
  wire [8:0] _T_334; // @[Shift.scala 91:22]
  wire [2:0] _T_335; // @[Shift.scala 92:77]
  wire [4:0] _T_336; // @[Shift.scala 90:30]
  wire [3:0] _T_337; // @[Shift.scala 90:48]
  wire  _T_338; // @[Shift.scala 90:57]
  wire [4:0] _GEN_20; // @[Shift.scala 90:39]
  wire [4:0] _T_339; // @[Shift.scala 90:39]
  wire  _T_340; // @[Shift.scala 12:21]
  wire  _T_341; // @[Shift.scala 12:21]
  wire [3:0] _T_343; // @[Bitwise.scala 71:12]
  wire [8:0] _T_344; // @[Cat.scala 29:58]
  wire [8:0] _T_345; // @[Shift.scala 91:22]
  wire [1:0] _T_346; // @[Shift.scala 92:77]
  wire [6:0] _T_347; // @[Shift.scala 90:30]
  wire [1:0] _T_348; // @[Shift.scala 90:48]
  wire  _T_349; // @[Shift.scala 90:57]
  wire [6:0] _GEN_21; // @[Shift.scala 90:39]
  wire [6:0] _T_350; // @[Shift.scala 90:39]
  wire  _T_351; // @[Shift.scala 12:21]
  wire  _T_352; // @[Shift.scala 12:21]
  wire [1:0] _T_354; // @[Bitwise.scala 71:12]
  wire [8:0] _T_355; // @[Cat.scala 29:58]
  wire [8:0] _T_356; // @[Shift.scala 91:22]
  wire  _T_357; // @[Shift.scala 92:77]
  wire [7:0] _T_358; // @[Shift.scala 90:30]
  wire  _T_359; // @[Shift.scala 90:48]
  wire [7:0] _GEN_22; // @[Shift.scala 90:39]
  wire [7:0] _T_361; // @[Shift.scala 90:39]
  wire  _T_363; // @[Shift.scala 12:21]
  wire [8:0] _T_364; // @[Cat.scala 29:58]
  wire [8:0] _T_365; // @[Shift.scala 91:22]
  wire [8:0] _T_368; // @[Bitwise.scala 71:12]
  wire [8:0] _T_369; // @[Shift.scala 39:10]
  wire  _T_370; // @[convert.scala 55:31]
  wire  _T_371; // @[convert.scala 56:31]
  wire  _T_372; // @[convert.scala 57:31]
  wire  _T_373; // @[convert.scala 58:31]
  wire [5:0] _T_374; // @[convert.scala 59:69]
  wire  _T_375; // @[convert.scala 59:81]
  wire  _T_376; // @[convert.scala 59:50]
  wire  _T_378; // @[convert.scala 60:81]
  wire  _T_379; // @[convert.scala 61:44]
  wire  _T_380; // @[convert.scala 61:52]
  wire  _T_381; // @[convert.scala 61:36]
  wire  _T_382; // @[convert.scala 62:63]
  wire  _T_383; // @[convert.scala 62:103]
  wire  _T_384; // @[convert.scala 62:60]
  wire [5:0] _GEN_23; // @[convert.scala 63:56]
  wire [5:0] _T_387; // @[convert.scala 63:56]
  wire [6:0] _T_388; // @[Cat.scala 29:58]
  wire [6:0] _T_390; // @[Mux.scala 87:16]
  assign _T_1 = io_A[6]; // @[convert.scala 18:24]
  assign _T_2 = io_A[5]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[5:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[4:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[4:1]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[3:2]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8 != 2'h0; // @[LZD.scala 39:14]
  assign _T_10 = _T_8[1]; // @[LZD.scala 39:21]
  assign _T_11 = _T_8[0]; // @[LZD.scala 39:30]
  assign _T_12 = ~ _T_11; // @[LZD.scala 39:27]
  assign _T_13 = _T_10 | _T_12; // @[LZD.scala 39:25]
  assign _T_14 = {_T_9,_T_13}; // @[Cat.scala 29:58]
  assign _T_15 = _T_7[1:0]; // @[LZD.scala 44:32]
  assign _T_16 = _T_15 != 2'h0; // @[LZD.scala 39:14]
  assign _T_17 = _T_15[1]; // @[LZD.scala 39:21]
  assign _T_18 = _T_15[0]; // @[LZD.scala 39:30]
  assign _T_19 = ~ _T_18; // @[LZD.scala 39:27]
  assign _T_20 = _T_17 | _T_19; // @[LZD.scala 39:25]
  assign _T_21 = {_T_16,_T_20}; // @[Cat.scala 29:58]
  assign _T_22 = _T_14[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22 | _T_23; // @[LZD.scala 49:16]
  assign _T_25 = ~ _T_23; // @[LZD.scala 49:27]
  assign _T_26 = _T_22 | _T_25; // @[LZD.scala 49:25]
  assign _T_27 = _T_14[0:0]; // @[LZD.scala 49:47]
  assign _T_28 = _T_21[0:0]; // @[LZD.scala 49:59]
  assign _T_29 = _T_22 ? _T_27 : _T_28; // @[LZD.scala 49:35]
  assign _T_31 = {_T_24,_T_26,_T_29}; // @[Cat.scala 29:58]
  assign _T_32 = _T_6[0:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_31[2]; // @[Shift.scala 12:21]
  assign _T_36 = {1'h1,_T_32}; // @[Cat.scala 29:58]
  assign _T_37 = _T_31[1:0]; // @[LZD.scala 55:32]
  assign _T_38 = _T_34 ? _T_37 : _T_36; // @[LZD.scala 55:20]
  assign _T_39 = {_T_34,_T_38}; // @[Cat.scala 29:58]
  assign _T_40 = ~ _T_39; // @[convert.scala 21:22]
  assign _T_41 = io_A[3:0]; // @[convert.scala 22:36]
  assign _T_42 = _T_40 < 3'h4; // @[Shift.scala 16:24]
  assign _T_43 = _T_40[1:0]; // @[Shift.scala 17:37]
  assign _T_44 = _T_43[1]; // @[Shift.scala 12:21]
  assign _T_45 = _T_41[1:0]; // @[Shift.scala 64:52]
  assign _T_47 = {_T_45,2'h0}; // @[Cat.scala 29:58]
  assign _T_48 = _T_44 ? _T_47 : _T_41; // @[Shift.scala 64:27]
  assign _T_49 = _T_43[0:0]; // @[Shift.scala 66:70]
  assign _T_51 = _T_48[2:0]; // @[Shift.scala 64:52]
  assign _T_52 = {_T_51,1'h0}; // @[Cat.scala 29:58]
  assign _T_53 = _T_49 ? _T_52 : _T_48; // @[Shift.scala 64:27]
  assign decA_fraction = _T_42 ? _T_53 : 4'h0; // @[Shift.scala 16:10]
  assign _T_57 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_59 = _T_3 ? _T_40 : _T_39; // @[convert.scala 25:42]
  assign _T_60 = {_T_57,_T_59}; // @[Cat.scala 29:58]
  assign _T_62 = io_A[5:0]; // @[convert.scala 29:56]
  assign _T_63 = _T_62 != 6'h0; // @[convert.scala 29:60]
  assign _T_64 = ~ _T_63; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_64; // @[convert.scala 29:39]
  assign _T_67 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_67 & _T_64; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_60); // @[convert.scala 32:24]
  assign _T_76 = io_B[6]; // @[convert.scala 18:24]
  assign _T_77 = io_B[5]; // @[convert.scala 18:40]
  assign _T_78 = _T_76 ^ _T_77; // @[convert.scala 18:36]
  assign _T_79 = io_B[5:1]; // @[convert.scala 19:24]
  assign _T_80 = io_B[4:0]; // @[convert.scala 19:43]
  assign _T_81 = _T_79 ^ _T_80; // @[convert.scala 19:39]
  assign _T_82 = _T_81[4:1]; // @[LZD.scala 43:32]
  assign _T_83 = _T_82[3:2]; // @[LZD.scala 43:32]
  assign _T_84 = _T_83 != 2'h0; // @[LZD.scala 39:14]
  assign _T_85 = _T_83[1]; // @[LZD.scala 39:21]
  assign _T_86 = _T_83[0]; // @[LZD.scala 39:30]
  assign _T_87 = ~ _T_86; // @[LZD.scala 39:27]
  assign _T_88 = _T_85 | _T_87; // @[LZD.scala 39:25]
  assign _T_89 = {_T_84,_T_88}; // @[Cat.scala 29:58]
  assign _T_90 = _T_82[1:0]; // @[LZD.scala 44:32]
  assign _T_91 = _T_90 != 2'h0; // @[LZD.scala 39:14]
  assign _T_92 = _T_90[1]; // @[LZD.scala 39:21]
  assign _T_93 = _T_90[0]; // @[LZD.scala 39:30]
  assign _T_94 = ~ _T_93; // @[LZD.scala 39:27]
  assign _T_95 = _T_92 | _T_94; // @[LZD.scala 39:25]
  assign _T_96 = {_T_91,_T_95}; // @[Cat.scala 29:58]
  assign _T_97 = _T_89[1]; // @[Shift.scala 12:21]
  assign _T_98 = _T_96[1]; // @[Shift.scala 12:21]
  assign _T_99 = _T_97 | _T_98; // @[LZD.scala 49:16]
  assign _T_100 = ~ _T_98; // @[LZD.scala 49:27]
  assign _T_101 = _T_97 | _T_100; // @[LZD.scala 49:25]
  assign _T_102 = _T_89[0:0]; // @[LZD.scala 49:47]
  assign _T_103 = _T_96[0:0]; // @[LZD.scala 49:59]
  assign _T_104 = _T_97 ? _T_102 : _T_103; // @[LZD.scala 49:35]
  assign _T_106 = {_T_99,_T_101,_T_104}; // @[Cat.scala 29:58]
  assign _T_107 = _T_81[0:0]; // @[LZD.scala 44:32]
  assign _T_109 = _T_106[2]; // @[Shift.scala 12:21]
  assign _T_111 = {1'h1,_T_107}; // @[Cat.scala 29:58]
  assign _T_112 = _T_106[1:0]; // @[LZD.scala 55:32]
  assign _T_113 = _T_109 ? _T_112 : _T_111; // @[LZD.scala 55:20]
  assign _T_114 = {_T_109,_T_113}; // @[Cat.scala 29:58]
  assign _T_115 = ~ _T_114; // @[convert.scala 21:22]
  assign _T_116 = io_B[3:0]; // @[convert.scala 22:36]
  assign _T_117 = _T_115 < 3'h4; // @[Shift.scala 16:24]
  assign _T_118 = _T_115[1:0]; // @[Shift.scala 17:37]
  assign _T_119 = _T_118[1]; // @[Shift.scala 12:21]
  assign _T_120 = _T_116[1:0]; // @[Shift.scala 64:52]
  assign _T_122 = {_T_120,2'h0}; // @[Cat.scala 29:58]
  assign _T_123 = _T_119 ? _T_122 : _T_116; // @[Shift.scala 64:27]
  assign _T_124 = _T_118[0:0]; // @[Shift.scala 66:70]
  assign _T_126 = _T_123[2:0]; // @[Shift.scala 64:52]
  assign _T_127 = {_T_126,1'h0}; // @[Cat.scala 29:58]
  assign _T_128 = _T_124 ? _T_127 : _T_123; // @[Shift.scala 64:27]
  assign decB_fraction = _T_117 ? _T_128 : 4'h0; // @[Shift.scala 16:10]
  assign _T_132 = _T_78 == 1'h0; // @[convert.scala 25:26]
  assign _T_134 = _T_78 ? _T_115 : _T_114; // @[convert.scala 25:42]
  assign _T_135 = {_T_132,_T_134}; // @[Cat.scala 29:58]
  assign _T_137 = io_B[5:0]; // @[convert.scala 29:56]
  assign _T_138 = _T_137 != 6'h0; // @[convert.scala 29:60]
  assign _T_139 = ~ _T_138; // @[convert.scala 29:41]
  assign decB_isNaR = _T_76 & _T_139; // @[convert.scala 29:39]
  assign _T_142 = _T_76 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_142 & _T_139; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_135); // @[convert.scala 32:24]
  assign _T_151 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_152 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_151,_T_152,decA_fraction,3'h0}; // @[Cat.scala 29:58]
  assign _T_155 = ~ _T_76; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_76,_T_155,decB_fraction,5'h0}; // @[Cat.scala 29:58]
  assign _T_158 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_158 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_159 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_160 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_161 = _T_160 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_162 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_163 = decA_isZero & _T_162; // @[PositDivisionSqrt.scala 94:43]
  assign _T_164 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_165 = _T_163 & _T_164; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_166 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_167 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_166 & _T_167; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_166 & _T_67; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_170 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_170; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 4'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_171 = sigX_Z[10]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_172 = sigX_Z[8]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_171 ^ _T_172; // @[PositDivisionSqrt.scala 113:50]
  assign _T_173 = cycleNum == 4'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_173 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_174 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_175 = _T_174 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_176 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_177 = entering & _T_176; // @[PositDivisionSqrt.scala 117:30]
  assign _T_179 = io_sqrtOp ? 4'h9 : 4'hb; // @[PositDivisionSqrt.scala 119:26]
  assign _T_180 = entering_normalCase ? _T_179 : 4'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{3'd0}, _T_177}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_181 = _GEN_9 | _T_180; // @[PositDivisionSqrt.scala 117:64]
  assign _T_183 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_184 = _T_174 & _T_183; // @[PositDivisionSqrt.scala 123:27]
  assign _T_186 = cycleNum - 4'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_187 = _T_184 ? _T_186 : 4'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _T_188 = _T_181 | _T_187; // @[PositDivisionSqrt.scala 122:64]
  assign _T_190 = _T_174 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_10 = {{3'd0}, _T_190}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_192 = _T_188 | _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  assign _T_193 = decA_scale[3:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_195 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_196 = entering_normalCase & _T_195; // @[PositDivisionSqrt.scala 137:28]
  assign _T_197 = 16'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign _T_198 = _T_197[15:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_199 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_200 = ready & _T_199; // @[PositDivisionSqrt.scala 148:23]
  assign _T_201 = _T_200 ? sigA_S : 11'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_202 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_203 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_204 = _T_203[10:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_205 = _T_202 ? _T_204 : 11'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_206 = _T_201 | _T_205; // @[PositDivisionSqrt.scala 148:66]
  assign _T_207 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_208 = _T_207 ? rem_Z : 11'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_206 | _T_208; // @[PositDivisionSqrt.scala 149:66]
  assign _T_210 = ready & _T_195; // @[PositDivisionSqrt.scala 152:29]
  assign _T_211 = _T_210 ? sigB_S : 11'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_212 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_213 = _T_212 ? 8'h80 : 8'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_11 = {{3'd0}, _T_213}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_214 = _T_211 | _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  assign _T_216 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_217 = _T_207 & _T_216; // @[PositDivisionSqrt.scala 154:30]
  assign _T_218 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_221 = {signB_Z,_T_218,fractB_Z,5'h0}; // @[Cat.scala 29:58]
  assign _T_222 = _T_217 ? _T_221 : 11'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_223 = _T_214 | _T_222; // @[PositDivisionSqrt.scala 153:93]
  assign _T_225 = _T_207 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_226 = rem[10:10]; // @[PositDivisionSqrt.scala 156:83]
  assign _T_228 = _T_226 ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign bitMask = _T_198[9:0]; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  assign _GEN_12 = {{3'd0}, _T_228}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_229 = bitMask & _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_13 = {{1'd0}, _T_229}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_230 = sigX_Z | _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  assign _T_231 = bitMask[9:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_14 = {{2'd0}, _T_231}; // @[PositDivisionSqrt.scala 156:89]
  assign _T_232 = _T_230 | _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  assign _T_233 = _T_225 ? _T_232 : 11'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_223 | _T_233; // @[PositDivisionSqrt.scala 154:93]
  assign _T_235 = trialTerm[10:10]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_236 = _T_226 ^ _T_235; // @[PositDivisionSqrt.scala 162:40]
  assign _T_239 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_241 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_242 = _T_236 ? _T_239 : _T_241; // @[PositDivisionSqrt.scala 161:92]
  assign _T_247 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_248 = _T_247[10:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_250 = _T_248 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_254 = _T_248 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_255 = _T_236 ? _T_250 : _T_254; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_242 : _T_255; // @[PositDivisionSqrt.scala 159:27]
  assign _T_256 = trialRem != 11'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_256 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_257 = rem != 11'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_257 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_259 = trialRem[10:10]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_260 = _T_235 ^ _T_259; // @[PositDivisionSqrt.scala 176:49]
  assign _T_261 = ~ _T_260; // @[PositDivisionSqrt.scala 176:29]
  assign _T_262 = sigX_Z[10:10]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_263 = ~ _T_262; // @[PositDivisionSqrt.scala 178:49]
  assign _T_265 = remIsZero ? _T_262 : _T_261; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_263 : _T_265; // @[Mux.scala 87:16]
  assign _T_266 = cycleNum > 4'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_267 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_268 = _T_266 & _T_267; // @[PositDivisionSqrt.scala 183:48]
  assign _T_269 = entering_normalCase | _T_268; // @[PositDivisionSqrt.scala 183:28]
  assign _T_272 = _T_207 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_273 = entering_normalCase | _T_272; // @[PositDivisionSqrt.scala 187:28]
  assign _T_276 = {newBit, 10'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_277 = _T_210 ? _T_276 : 11'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_279 = _T_212 ? 9'h100 : 9'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_15 = {{2'd0}, _T_279}; // @[PositDivisionSqrt.scala 188:78]
  assign _T_280 = _T_277 | _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  assign _GEN_16 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_282 = sigX_Z | _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  assign _T_283 = _T_207 ? _T_282 : 11'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_284 = _T_280 | _T_283; // @[PositDivisionSqrt.scala 189:78]
  assign _T_286 = {_T_262, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_286 : {{1'd0}, _T_262}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_17 = {{9'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  assign _T_289 = realSigX[7:4]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_290 = realSigX[6:3]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_289 : _T_290; // @[PositDivisionSqrt.scala 198:21]
  assign _T_291 = realSigX[10]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_292 = realSigX[8]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_293 = _T_291 ^ _T_292; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_293; // @[PositDivisionSqrt.scala 205:23]
  assign _T_295 = realSigX[7]; // @[PositDivisionSqrt.scala 206:56]
  assign notNeedSubTwo = _T_291 ^ _T_295; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_296 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_296; // @[PositDivisionSqrt.scala 208:36]
  assign _T_297 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_298 = {1'b0,$signed(_T_297)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_18 = {{2{_T_298[2]}},_T_298}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_300 = $signed(scale_Z) - $signed(_GEN_18); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_300); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-5'sh6); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(5'sh5); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[10:10]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_302 = underflow ? $signed(-5'sh6) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_303 = overflow ? $signed(5'sh5) : $signed(_T_302); // @[Mux.scala 87:16]
  assign _T_304 = realSigX[3:1]; // @[PositDivisionSqrt.scala 224:48]
  assign _T_305 = realSigX[2:0]; // @[PositDivisionSqrt.scala 224:64]
  assign decQ_grs = scaleNotChange ? _T_304 : _T_305; // @[PositDivisionSqrt.scala 224:23]
  assign outValid = cycleNum == 4'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_19 = _T_303[3:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_19); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_312 = decQ_scale[3:3]; // @[convert.scala 49:36]
  assign _T_314 = ~ decQ_scale; // @[convert.scala 50:36]
  assign _T_315 = $signed(_T_314); // @[convert.scala 50:36]
  assign _T_316 = _T_312 ? $signed(_T_315) : $signed(decQ_scale); // @[convert.scala 50:28]
  assign _T_317 = _T_312 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_318 = ~ _T_317; // @[convert.scala 53:34]
  assign _T_321 = {_T_318,_T_317,realFrac,decQ_grs}; // @[Cat.scala 29:58]
  assign _T_322 = $unsigned(_T_316); // @[Shift.scala 39:17]
  assign _T_323 = _T_322 < 4'h9; // @[Shift.scala 39:24]
  assign _T_325 = _T_321[8:8]; // @[Shift.scala 90:30]
  assign _T_326 = _T_321[7:0]; // @[Shift.scala 90:48]
  assign _T_327 = _T_326 != 8'h0; // @[Shift.scala 90:57]
  assign _T_328 = _T_325 | _T_327; // @[Shift.scala 90:39]
  assign _T_329 = _T_322[3]; // @[Shift.scala 12:21]
  assign _T_330 = _T_321[8]; // @[Shift.scala 12:21]
  assign _T_332 = _T_330 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_333 = {_T_332,_T_328}; // @[Cat.scala 29:58]
  assign _T_334 = _T_329 ? _T_333 : _T_321; // @[Shift.scala 91:22]
  assign _T_335 = _T_322[2:0]; // @[Shift.scala 92:77]
  assign _T_336 = _T_334[8:4]; // @[Shift.scala 90:30]
  assign _T_337 = _T_334[3:0]; // @[Shift.scala 90:48]
  assign _T_338 = _T_337 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{4'd0}, _T_338}; // @[Shift.scala 90:39]
  assign _T_339 = _T_336 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_340 = _T_335[2]; // @[Shift.scala 12:21]
  assign _T_341 = _T_334[8]; // @[Shift.scala 12:21]
  assign _T_343 = _T_341 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_344 = {_T_343,_T_339}; // @[Cat.scala 29:58]
  assign _T_345 = _T_340 ? _T_344 : _T_334; // @[Shift.scala 91:22]
  assign _T_346 = _T_335[1:0]; // @[Shift.scala 92:77]
  assign _T_347 = _T_345[8:2]; // @[Shift.scala 90:30]
  assign _T_348 = _T_345[1:0]; // @[Shift.scala 90:48]
  assign _T_349 = _T_348 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{6'd0}, _T_349}; // @[Shift.scala 90:39]
  assign _T_350 = _T_347 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_351 = _T_346[1]; // @[Shift.scala 12:21]
  assign _T_352 = _T_345[8]; // @[Shift.scala 12:21]
  assign _T_354 = _T_352 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_355 = {_T_354,_T_350}; // @[Cat.scala 29:58]
  assign _T_356 = _T_351 ? _T_355 : _T_345; // @[Shift.scala 91:22]
  assign _T_357 = _T_346[0:0]; // @[Shift.scala 92:77]
  assign _T_358 = _T_356[8:1]; // @[Shift.scala 90:30]
  assign _T_359 = _T_356[0:0]; // @[Shift.scala 90:48]
  assign _GEN_22 = {{7'd0}, _T_359}; // @[Shift.scala 90:39]
  assign _T_361 = _T_358 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_363 = _T_356[8]; // @[Shift.scala 12:21]
  assign _T_364 = {_T_363,_T_361}; // @[Cat.scala 29:58]
  assign _T_365 = _T_357 ? _T_364 : _T_356; // @[Shift.scala 91:22]
  assign _T_368 = _T_330 ? 9'h1ff : 9'h0; // @[Bitwise.scala 71:12]
  assign _T_369 = _T_323 ? _T_365 : _T_368; // @[Shift.scala 39:10]
  assign _T_370 = _T_369[3]; // @[convert.scala 55:31]
  assign _T_371 = _T_369[2]; // @[convert.scala 56:31]
  assign _T_372 = _T_369[1]; // @[convert.scala 57:31]
  assign _T_373 = _T_369[0]; // @[convert.scala 58:31]
  assign _T_374 = _T_369[8:3]; // @[convert.scala 59:69]
  assign _T_375 = _T_374 != 6'h0; // @[convert.scala 59:81]
  assign _T_376 = ~ _T_375; // @[convert.scala 59:50]
  assign _T_378 = _T_374 == 6'h3f; // @[convert.scala 60:81]
  assign _T_379 = _T_370 | _T_372; // @[convert.scala 61:44]
  assign _T_380 = _T_379 | _T_373; // @[convert.scala 61:52]
  assign _T_381 = _T_371 & _T_380; // @[convert.scala 61:36]
  assign _T_382 = ~ _T_378; // @[convert.scala 62:63]
  assign _T_383 = _T_382 & _T_381; // @[convert.scala 62:103]
  assign _T_384 = _T_376 | _T_383; // @[convert.scala 62:60]
  assign _GEN_23 = {{5'd0}, _T_384}; // @[convert.scala 63:56]
  assign _T_387 = _T_374 + _GEN_23; // @[convert.scala 63:56]
  assign _T_388 = {decQ_sign,_T_387}; // @[Cat.scala 29:58]
  assign _T_390 = isZero_Z ? 7'h0 : _T_388; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_216; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 7'h40 : _T_390; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[10:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 4'h0;
    end else begin
      if (_T_175) begin
        cycleNum <= _T_192;
      end
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_159;
      end else begin
        isNaR_Z <= _T_161;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_165;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_193[2]}},_T_193};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_196) begin
      signB_Z <= _T_76;
    end
    if (_T_196) begin
      if (_T_117) begin
        if (_T_124) begin
          fractB_Z <= _T_127;
        end else begin
          if (_T_119) begin
            fractB_Z <= _T_122;
          end else begin
            fractB_Z <= _T_116;
          end
        end
      end else begin
        fractB_Z <= 4'h0;
      end
    end
    if (_T_269) begin
      if (ready) begin
        if (_T_236) begin
          rem_Z <= _T_239;
        end else begin
          rem_Z <= _T_241;
        end
      end else begin
        if (_T_236) begin
          rem_Z <= _T_250;
        end else begin
          rem_Z <= _T_254;
        end
      end
    end
    if (_T_273) begin
      sigX_Z <= _T_284;
    end
  end
endmodule
