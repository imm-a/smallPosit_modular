module FMAEnc8_2(
  input        clock,
  input        reset,
  input        io_inValid_phase2,
  input  [9:0] io_signSumSig,
  input        io_sumSign,
  input  [5:0] io_greaterScale,
  input        io_outIsNaR_phase2,
  output [7:0] io_F,
  output       io_outValid
);
  wire [8:0] _T; // @[FMAEnc.scala 35:36]
  wire [8:0] _T_1; // @[FMAEnc.scala 35:74]
  wire [8:0] sumXor; // @[FMAEnc.scala 35:54]
  wire [7:0] _T_2; // @[LZD.scala 43:32]
  wire [3:0] _T_3; // @[LZD.scala 43:32]
  wire [1:0] _T_4; // @[LZD.scala 43:32]
  wire  _T_5; // @[LZD.scala 39:14]
  wire  _T_6; // @[LZD.scala 39:21]
  wire  _T_7; // @[LZD.scala 39:30]
  wire  _T_8; // @[LZD.scala 39:27]
  wire  _T_9; // @[LZD.scala 39:25]
  wire [1:0] _T_10; // @[Cat.scala 29:58]
  wire [1:0] _T_11; // @[LZD.scala 44:32]
  wire  _T_12; // @[LZD.scala 39:14]
  wire  _T_13; // @[LZD.scala 39:21]
  wire  _T_14; // @[LZD.scala 39:30]
  wire  _T_15; // @[LZD.scala 39:27]
  wire  _T_16; // @[LZD.scala 39:25]
  wire [1:0] _T_17; // @[Cat.scala 29:58]
  wire  _T_18; // @[Shift.scala 12:21]
  wire  _T_19; // @[Shift.scala 12:21]
  wire  _T_20; // @[LZD.scala 49:16]
  wire  _T_21; // @[LZD.scala 49:27]
  wire  _T_22; // @[LZD.scala 49:25]
  wire  _T_23; // @[LZD.scala 49:47]
  wire  _T_24; // @[LZD.scala 49:59]
  wire  _T_25; // @[LZD.scala 49:35]
  wire [2:0] _T_27; // @[Cat.scala 29:58]
  wire [3:0] _T_28; // @[LZD.scala 44:32]
  wire [1:0] _T_29; // @[LZD.scala 43:32]
  wire  _T_30; // @[LZD.scala 39:14]
  wire  _T_31; // @[LZD.scala 39:21]
  wire  _T_32; // @[LZD.scala 39:30]
  wire  _T_33; // @[LZD.scala 39:27]
  wire  _T_34; // @[LZD.scala 39:25]
  wire [1:0] _T_35; // @[Cat.scala 29:58]
  wire [1:0] _T_36; // @[LZD.scala 44:32]
  wire  _T_37; // @[LZD.scala 39:14]
  wire  _T_38; // @[LZD.scala 39:21]
  wire  _T_39; // @[LZD.scala 39:30]
  wire  _T_40; // @[LZD.scala 39:27]
  wire  _T_41; // @[LZD.scala 39:25]
  wire [1:0] _T_42; // @[Cat.scala 29:58]
  wire  _T_43; // @[Shift.scala 12:21]
  wire  _T_44; // @[Shift.scala 12:21]
  wire  _T_45; // @[LZD.scala 49:16]
  wire  _T_46; // @[LZD.scala 49:27]
  wire  _T_47; // @[LZD.scala 49:25]
  wire  _T_48; // @[LZD.scala 49:47]
  wire  _T_49; // @[LZD.scala 49:59]
  wire  _T_50; // @[LZD.scala 49:35]
  wire [2:0] _T_52; // @[Cat.scala 29:58]
  wire  _T_53; // @[Shift.scala 12:21]
  wire  _T_54; // @[Shift.scala 12:21]
  wire  _T_55; // @[LZD.scala 49:16]
  wire  _T_56; // @[LZD.scala 49:27]
  wire  _T_57; // @[LZD.scala 49:25]
  wire [1:0] _T_58; // @[LZD.scala 49:47]
  wire [1:0] _T_59; // @[LZD.scala 49:59]
  wire [1:0] _T_60; // @[LZD.scala 49:35]
  wire [3:0] _T_62; // @[Cat.scala 29:58]
  wire  _T_63; // @[LZD.scala 44:32]
  wire  _T_65; // @[Shift.scala 12:21]
  wire [2:0] _T_68; // @[Cat.scala 29:58]
  wire [2:0] _T_69; // @[LZD.scala 55:32]
  wire [2:0] _T_70; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [3:0] shiftValue; // @[FMAEnc.scala 37:24]
  wire [7:0] _T_71; // @[FMAEnc.scala 38:41]
  wire  _T_72; // @[Shift.scala 16:24]
  wire [2:0] _T_73; // @[Shift.scala 17:37]
  wire  _T_74; // @[Shift.scala 12:21]
  wire [3:0] _T_75; // @[Shift.scala 64:52]
  wire [7:0] _T_77; // @[Cat.scala 29:58]
  wire [7:0] _T_78; // @[Shift.scala 64:27]
  wire [1:0] _T_79; // @[Shift.scala 66:70]
  wire  _T_80; // @[Shift.scala 12:21]
  wire [5:0] _T_81; // @[Shift.scala 64:52]
  wire [7:0] _T_83; // @[Cat.scala 29:58]
  wire [7:0] _T_84; // @[Shift.scala 64:27]
  wire  _T_85; // @[Shift.scala 66:70]
  wire [6:0] _T_87; // @[Shift.scala 64:52]
  wire [7:0] _T_88; // @[Cat.scala 29:58]
  wire [7:0] _T_89; // @[Shift.scala 64:27]
  wire [7:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [5:0] _T_91; // @[FMAEnc.scala 41:39]
  wire [5:0] _T_92; // @[FMAEnc.scala 41:39]
  wire [4:0] _T_93; // @[Cat.scala 29:58]
  wire [4:0] _T_94; // @[FMAEnc.scala 41:64]
  wire [5:0] _GEN_2; // @[FMAEnc.scala 41:45]
  wire [5:0] _T_96; // @[FMAEnc.scala 41:45]
  wire [5:0] sumScale; // @[FMAEnc.scala 41:45]
  wire [2:0] sumFrac; // @[FMAEnc.scala 42:41]
  wire [4:0] grsTmp; // @[FMAEnc.scala 45:41]
  wire [1:0] _T_97; // @[FMAEnc.scala 48:40]
  wire [2:0] _T_98; // @[FMAEnc.scala 48:56]
  wire  _T_99; // @[FMAEnc.scala 48:60]
  wire  underflow; // @[FMAEnc.scala 55:32]
  wire  overflow; // @[FMAEnc.scala 56:32]
  wire  _T_100; // @[FMAEnc.scala 65:35]
  wire  decF_isZero; // @[FMAEnc.scala 65:20]
  wire [5:0] _T_102; // @[Mux.scala 87:16]
  wire [5:0] decF_scale; // @[Mux.scala 87:16]
  wire [1:0] _T_104; // @[convert.scala 46:61]
  wire [1:0] _T_105; // @[convert.scala 46:52]
  wire [1:0] _T_107; // @[convert.scala 46:42]
  wire [3:0] _T_108; // @[convert.scala 48:34]
  wire  _T_109; // @[convert.scala 49:36]
  wire [3:0] _T_111; // @[convert.scala 50:36]
  wire [3:0] _T_112; // @[convert.scala 50:36]
  wire [3:0] _T_113; // @[convert.scala 50:28]
  wire  _T_114; // @[convert.scala 51:31]
  wire  _T_115; // @[convert.scala 52:43]
  wire [9:0] _T_119; // @[Cat.scala 29:58]
  wire [3:0] _T_120; // @[Shift.scala 39:17]
  wire  _T_121; // @[Shift.scala 39:24]
  wire [1:0] _T_123; // @[Shift.scala 90:30]
  wire [7:0] _T_124; // @[Shift.scala 90:48]
  wire  _T_125; // @[Shift.scala 90:57]
  wire [1:0] _GEN_3; // @[Shift.scala 90:39]
  wire [1:0] _T_126; // @[Shift.scala 90:39]
  wire  _T_127; // @[Shift.scala 12:21]
  wire  _T_128; // @[Shift.scala 12:21]
  wire [7:0] _T_130; // @[Bitwise.scala 71:12]
  wire [9:0] _T_131; // @[Cat.scala 29:58]
  wire [9:0] _T_132; // @[Shift.scala 91:22]
  wire [2:0] _T_133; // @[Shift.scala 92:77]
  wire [5:0] _T_134; // @[Shift.scala 90:30]
  wire [3:0] _T_135; // @[Shift.scala 90:48]
  wire  _T_136; // @[Shift.scala 90:57]
  wire [5:0] _GEN_4; // @[Shift.scala 90:39]
  wire [5:0] _T_137; // @[Shift.scala 90:39]
  wire  _T_138; // @[Shift.scala 12:21]
  wire  _T_139; // @[Shift.scala 12:21]
  wire [3:0] _T_141; // @[Bitwise.scala 71:12]
  wire [9:0] _T_142; // @[Cat.scala 29:58]
  wire [9:0] _T_143; // @[Shift.scala 91:22]
  wire [1:0] _T_144; // @[Shift.scala 92:77]
  wire [7:0] _T_145; // @[Shift.scala 90:30]
  wire [1:0] _T_146; // @[Shift.scala 90:48]
  wire  _T_147; // @[Shift.scala 90:57]
  wire [7:0] _GEN_5; // @[Shift.scala 90:39]
  wire [7:0] _T_148; // @[Shift.scala 90:39]
  wire  _T_149; // @[Shift.scala 12:21]
  wire  _T_150; // @[Shift.scala 12:21]
  wire [1:0] _T_152; // @[Bitwise.scala 71:12]
  wire [9:0] _T_153; // @[Cat.scala 29:58]
  wire [9:0] _T_154; // @[Shift.scala 91:22]
  wire  _T_155; // @[Shift.scala 92:77]
  wire [8:0] _T_156; // @[Shift.scala 90:30]
  wire  _T_157; // @[Shift.scala 90:48]
  wire [8:0] _GEN_6; // @[Shift.scala 90:39]
  wire [8:0] _T_159; // @[Shift.scala 90:39]
  wire  _T_161; // @[Shift.scala 12:21]
  wire [9:0] _T_162; // @[Cat.scala 29:58]
  wire [9:0] _T_163; // @[Shift.scala 91:22]
  wire [9:0] _T_166; // @[Bitwise.scala 71:12]
  wire [9:0] _T_167; // @[Shift.scala 39:10]
  wire  _T_168; // @[convert.scala 55:31]
  wire  _T_169; // @[convert.scala 56:31]
  wire  _T_170; // @[convert.scala 57:31]
  wire  _T_171; // @[convert.scala 58:31]
  wire [6:0] _T_172; // @[convert.scala 59:69]
  wire  _T_173; // @[convert.scala 59:81]
  wire  _T_174; // @[convert.scala 59:50]
  wire  _T_176; // @[convert.scala 60:81]
  wire  _T_177; // @[convert.scala 61:44]
  wire  _T_178; // @[convert.scala 61:52]
  wire  _T_179; // @[convert.scala 61:36]
  wire  _T_180; // @[convert.scala 62:63]
  wire  _T_181; // @[convert.scala 62:103]
  wire  _T_182; // @[convert.scala 62:60]
  wire [6:0] _GEN_7; // @[convert.scala 63:56]
  wire [6:0] _T_185; // @[convert.scala 63:56]
  wire [7:0] _T_186; // @[Cat.scala 29:58]
  reg  _T_190; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [7:0] _T_194; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  assign _T = io_signSumSig[9:1]; // @[FMAEnc.scala 35:36]
  assign _T_1 = io_signSumSig[8:0]; // @[FMAEnc.scala 35:74]
  assign sumXor = _T ^ _T_1; // @[FMAEnc.scala 35:54]
  assign _T_2 = sumXor[8:1]; // @[LZD.scala 43:32]
  assign _T_3 = _T_2[7:4]; // @[LZD.scala 43:32]
  assign _T_4 = _T_3[3:2]; // @[LZD.scala 43:32]
  assign _T_5 = _T_4 != 2'h0; // @[LZD.scala 39:14]
  assign _T_6 = _T_4[1]; // @[LZD.scala 39:21]
  assign _T_7 = _T_4[0]; // @[LZD.scala 39:30]
  assign _T_8 = ~ _T_7; // @[LZD.scala 39:27]
  assign _T_9 = _T_6 | _T_8; // @[LZD.scala 39:25]
  assign _T_10 = {_T_5,_T_9}; // @[Cat.scala 29:58]
  assign _T_11 = _T_3[1:0]; // @[LZD.scala 44:32]
  assign _T_12 = _T_11 != 2'h0; // @[LZD.scala 39:14]
  assign _T_13 = _T_11[1]; // @[LZD.scala 39:21]
  assign _T_14 = _T_11[0]; // @[LZD.scala 39:30]
  assign _T_15 = ~ _T_14; // @[LZD.scala 39:27]
  assign _T_16 = _T_13 | _T_15; // @[LZD.scala 39:25]
  assign _T_17 = {_T_12,_T_16}; // @[Cat.scala 29:58]
  assign _T_18 = _T_10[1]; // @[Shift.scala 12:21]
  assign _T_19 = _T_17[1]; // @[Shift.scala 12:21]
  assign _T_20 = _T_18 | _T_19; // @[LZD.scala 49:16]
  assign _T_21 = ~ _T_19; // @[LZD.scala 49:27]
  assign _T_22 = _T_18 | _T_21; // @[LZD.scala 49:25]
  assign _T_23 = _T_10[0:0]; // @[LZD.scala 49:47]
  assign _T_24 = _T_17[0:0]; // @[LZD.scala 49:59]
  assign _T_25 = _T_18 ? _T_23 : _T_24; // @[LZD.scala 49:35]
  assign _T_27 = {_T_20,_T_22,_T_25}; // @[Cat.scala 29:58]
  assign _T_28 = _T_2[3:0]; // @[LZD.scala 44:32]
  assign _T_29 = _T_28[3:2]; // @[LZD.scala 43:32]
  assign _T_30 = _T_29 != 2'h0; // @[LZD.scala 39:14]
  assign _T_31 = _T_29[1]; // @[LZD.scala 39:21]
  assign _T_32 = _T_29[0]; // @[LZD.scala 39:30]
  assign _T_33 = ~ _T_32; // @[LZD.scala 39:27]
  assign _T_34 = _T_31 | _T_33; // @[LZD.scala 39:25]
  assign _T_35 = {_T_30,_T_34}; // @[Cat.scala 29:58]
  assign _T_36 = _T_28[1:0]; // @[LZD.scala 44:32]
  assign _T_37 = _T_36 != 2'h0; // @[LZD.scala 39:14]
  assign _T_38 = _T_36[1]; // @[LZD.scala 39:21]
  assign _T_39 = _T_36[0]; // @[LZD.scala 39:30]
  assign _T_40 = ~ _T_39; // @[LZD.scala 39:27]
  assign _T_41 = _T_38 | _T_40; // @[LZD.scala 39:25]
  assign _T_42 = {_T_37,_T_41}; // @[Cat.scala 29:58]
  assign _T_43 = _T_35[1]; // @[Shift.scala 12:21]
  assign _T_44 = _T_42[1]; // @[Shift.scala 12:21]
  assign _T_45 = _T_43 | _T_44; // @[LZD.scala 49:16]
  assign _T_46 = ~ _T_44; // @[LZD.scala 49:27]
  assign _T_47 = _T_43 | _T_46; // @[LZD.scala 49:25]
  assign _T_48 = _T_35[0:0]; // @[LZD.scala 49:47]
  assign _T_49 = _T_42[0:0]; // @[LZD.scala 49:59]
  assign _T_50 = _T_43 ? _T_48 : _T_49; // @[LZD.scala 49:35]
  assign _T_52 = {_T_45,_T_47,_T_50}; // @[Cat.scala 29:58]
  assign _T_53 = _T_27[2]; // @[Shift.scala 12:21]
  assign _T_54 = _T_52[2]; // @[Shift.scala 12:21]
  assign _T_55 = _T_53 | _T_54; // @[LZD.scala 49:16]
  assign _T_56 = ~ _T_54; // @[LZD.scala 49:27]
  assign _T_57 = _T_53 | _T_56; // @[LZD.scala 49:25]
  assign _T_58 = _T_27[1:0]; // @[LZD.scala 49:47]
  assign _T_59 = _T_52[1:0]; // @[LZD.scala 49:59]
  assign _T_60 = _T_53 ? _T_58 : _T_59; // @[LZD.scala 49:35]
  assign _T_62 = {_T_55,_T_57,_T_60}; // @[Cat.scala 29:58]
  assign _T_63 = sumXor[0:0]; // @[LZD.scala 44:32]
  assign _T_65 = _T_62[3]; // @[Shift.scala 12:21]
  assign _T_68 = {2'h3,_T_63}; // @[Cat.scala 29:58]
  assign _T_69 = _T_62[2:0]; // @[LZD.scala 55:32]
  assign _T_70 = _T_65 ? _T_69 : _T_68; // @[LZD.scala 55:20]
  assign sumLZD = {_T_65,_T_70}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[FMAEnc.scala 37:24]
  assign _T_71 = io_signSumSig[7:0]; // @[FMAEnc.scala 38:41]
  assign _T_72 = shiftValue < 4'h8; // @[Shift.scala 16:24]
  assign _T_73 = shiftValue[2:0]; // @[Shift.scala 17:37]
  assign _T_74 = _T_73[2]; // @[Shift.scala 12:21]
  assign _T_75 = _T_71[3:0]; // @[Shift.scala 64:52]
  assign _T_77 = {_T_75,4'h0}; // @[Cat.scala 29:58]
  assign _T_78 = _T_74 ? _T_77 : _T_71; // @[Shift.scala 64:27]
  assign _T_79 = _T_73[1:0]; // @[Shift.scala 66:70]
  assign _T_80 = _T_79[1]; // @[Shift.scala 12:21]
  assign _T_81 = _T_78[5:0]; // @[Shift.scala 64:52]
  assign _T_83 = {_T_81,2'h0}; // @[Cat.scala 29:58]
  assign _T_84 = _T_80 ? _T_83 : _T_78; // @[Shift.scala 64:27]
  assign _T_85 = _T_79[0:0]; // @[Shift.scala 66:70]
  assign _T_87 = _T_84[6:0]; // @[Shift.scala 64:52]
  assign _T_88 = {_T_87,1'h0}; // @[Cat.scala 29:58]
  assign _T_89 = _T_85 ? _T_88 : _T_84; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_72 ? _T_89 : 8'h0; // @[Shift.scala 16:10]
  assign _T_91 = $signed(io_greaterScale) + $signed(6'sh2); // @[FMAEnc.scala 41:39]
  assign _T_92 = $signed(_T_91); // @[FMAEnc.scala 41:39]
  assign _T_93 = {1'h1,_T_65,_T_70}; // @[Cat.scala 29:58]
  assign _T_94 = $signed(_T_93); // @[FMAEnc.scala 41:64]
  assign _GEN_2 = {{1{_T_94[4]}},_T_94}; // @[FMAEnc.scala 41:45]
  assign _T_96 = $signed(_T_92) + $signed(_GEN_2); // @[FMAEnc.scala 41:45]
  assign sumScale = $signed(_T_96); // @[FMAEnc.scala 41:45]
  assign sumFrac = normalFracTmp[7:5]; // @[FMAEnc.scala 42:41]
  assign grsTmp = normalFracTmp[4:0]; // @[FMAEnc.scala 45:41]
  assign _T_97 = grsTmp[4:3]; // @[FMAEnc.scala 48:40]
  assign _T_98 = grsTmp[2:0]; // @[FMAEnc.scala 48:56]
  assign _T_99 = _T_98 != 3'h0; // @[FMAEnc.scala 48:60]
  assign underflow = $signed(sumScale) < $signed(-6'sh19); // @[FMAEnc.scala 55:32]
  assign overflow = $signed(sumScale) > $signed(6'sh18); // @[FMAEnc.scala 56:32]
  assign _T_100 = io_signSumSig != 10'h0; // @[FMAEnc.scala 65:35]
  assign decF_isZero = ~ _T_100; // @[FMAEnc.scala 65:20]
  assign _T_102 = underflow ? $signed(-6'sh19) : $signed(sumScale); // @[Mux.scala 87:16]
  assign decF_scale = overflow ? $signed(6'sh18) : $signed(_T_102); // @[Mux.scala 87:16]
  assign _T_104 = decF_scale[1:0]; // @[convert.scala 46:61]
  assign _T_105 = ~ _T_104; // @[convert.scala 46:52]
  assign _T_107 = io_sumSign ? _T_105 : _T_104; // @[convert.scala 46:42]
  assign _T_108 = decF_scale[5:2]; // @[convert.scala 48:34]
  assign _T_109 = _T_108[3:3]; // @[convert.scala 49:36]
  assign _T_111 = ~ _T_108; // @[convert.scala 50:36]
  assign _T_112 = $signed(_T_111); // @[convert.scala 50:36]
  assign _T_113 = _T_109 ? $signed(_T_112) : $signed(_T_108); // @[convert.scala 50:28]
  assign _T_114 = _T_109 ^ io_sumSign; // @[convert.scala 51:31]
  assign _T_115 = ~ _T_114; // @[convert.scala 52:43]
  assign _T_119 = {_T_115,_T_114,_T_107,sumFrac,_T_97,_T_99}; // @[Cat.scala 29:58]
  assign _T_120 = $unsigned(_T_113); // @[Shift.scala 39:17]
  assign _T_121 = _T_120 < 4'ha; // @[Shift.scala 39:24]
  assign _T_123 = _T_119[9:8]; // @[Shift.scala 90:30]
  assign _T_124 = _T_119[7:0]; // @[Shift.scala 90:48]
  assign _T_125 = _T_124 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_3 = {{1'd0}, _T_125}; // @[Shift.scala 90:39]
  assign _T_126 = _T_123 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_127 = _T_120[3]; // @[Shift.scala 12:21]
  assign _T_128 = _T_119[9]; // @[Shift.scala 12:21]
  assign _T_130 = _T_128 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_131 = {_T_130,_T_126}; // @[Cat.scala 29:58]
  assign _T_132 = _T_127 ? _T_131 : _T_119; // @[Shift.scala 91:22]
  assign _T_133 = _T_120[2:0]; // @[Shift.scala 92:77]
  assign _T_134 = _T_132[9:4]; // @[Shift.scala 90:30]
  assign _T_135 = _T_132[3:0]; // @[Shift.scala 90:48]
  assign _T_136 = _T_135 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_4 = {{5'd0}, _T_136}; // @[Shift.scala 90:39]
  assign _T_137 = _T_134 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_138 = _T_133[2]; // @[Shift.scala 12:21]
  assign _T_139 = _T_132[9]; // @[Shift.scala 12:21]
  assign _T_141 = _T_139 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_142 = {_T_141,_T_137}; // @[Cat.scala 29:58]
  assign _T_143 = _T_138 ? _T_142 : _T_132; // @[Shift.scala 91:22]
  assign _T_144 = _T_133[1:0]; // @[Shift.scala 92:77]
  assign _T_145 = _T_143[9:2]; // @[Shift.scala 90:30]
  assign _T_146 = _T_143[1:0]; // @[Shift.scala 90:48]
  assign _T_147 = _T_146 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{7'd0}, _T_147}; // @[Shift.scala 90:39]
  assign _T_148 = _T_145 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_149 = _T_144[1]; // @[Shift.scala 12:21]
  assign _T_150 = _T_143[9]; // @[Shift.scala 12:21]
  assign _T_152 = _T_150 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_153 = {_T_152,_T_148}; // @[Cat.scala 29:58]
  assign _T_154 = _T_149 ? _T_153 : _T_143; // @[Shift.scala 91:22]
  assign _T_155 = _T_144[0:0]; // @[Shift.scala 92:77]
  assign _T_156 = _T_154[9:1]; // @[Shift.scala 90:30]
  assign _T_157 = _T_154[0:0]; // @[Shift.scala 90:48]
  assign _GEN_6 = {{8'd0}, _T_157}; // @[Shift.scala 90:39]
  assign _T_159 = _T_156 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_161 = _T_154[9]; // @[Shift.scala 12:21]
  assign _T_162 = {_T_161,_T_159}; // @[Cat.scala 29:58]
  assign _T_163 = _T_155 ? _T_162 : _T_154; // @[Shift.scala 91:22]
  assign _T_166 = _T_128 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_167 = _T_121 ? _T_163 : _T_166; // @[Shift.scala 39:10]
  assign _T_168 = _T_167[3]; // @[convert.scala 55:31]
  assign _T_169 = _T_167[2]; // @[convert.scala 56:31]
  assign _T_170 = _T_167[1]; // @[convert.scala 57:31]
  assign _T_171 = _T_167[0]; // @[convert.scala 58:31]
  assign _T_172 = _T_167[9:3]; // @[convert.scala 59:69]
  assign _T_173 = _T_172 != 7'h0; // @[convert.scala 59:81]
  assign _T_174 = ~ _T_173; // @[convert.scala 59:50]
  assign _T_176 = _T_172 == 7'h7f; // @[convert.scala 60:81]
  assign _T_177 = _T_168 | _T_170; // @[convert.scala 61:44]
  assign _T_178 = _T_177 | _T_171; // @[convert.scala 61:52]
  assign _T_179 = _T_169 & _T_178; // @[convert.scala 61:36]
  assign _T_180 = ~ _T_176; // @[convert.scala 62:63]
  assign _T_181 = _T_180 & _T_179; // @[convert.scala 62:103]
  assign _T_182 = _T_174 | _T_181; // @[convert.scala 62:60]
  assign _GEN_7 = {{6'd0}, _T_182}; // @[convert.scala 63:56]
  assign _T_185 = _T_172 + _GEN_7; // @[convert.scala 63:56]
  assign _T_186 = {io_sumSign,_T_185}; // @[Cat.scala 29:58]
  assign io_F = _T_194; // @[FMAEnc.scala 85:15]
  assign io_outValid = _T_190; // @[FMAEnc.scala 84:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_190 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_194 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_190 <= 1'h0;
    end else begin
      _T_190 <= io_inValid_phase2;
    end
    if (io_inValid_phase2) begin
      if (io_outIsNaR_phase2) begin
        _T_194 <= 8'h80;
      end else begin
        if (decF_isZero) begin
          _T_194 <= 8'h0;
        end else begin
          _T_194 <= _T_186;
        end
      end
    end
  end
endmodule
