module PositDivSqrter5_1(
  input        clock,
  input        reset,
  output       io_inReady,
  input        io_inValid,
  input        io_sqrtOp,
  input  [4:0] io_A,
  input  [4:0] io_B,
  output       io_diviValid,
  output       io_sqrtValid,
  output       io_invalidExc,
  output [4:0] io_Q
);
  reg [2:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [4:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg  fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [7:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [7:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [2:0] _T_4; // @[convert.scala 19:24]
  wire [2:0] _T_5; // @[convert.scala 19:43]
  wire [2:0] _T_6; // @[convert.scala 19:39]
  wire [1:0] _T_7; // @[LZD.scala 43:32]
  wire  _T_8; // @[LZD.scala 39:14]
  wire  _T_9; // @[LZD.scala 39:21]
  wire  _T_10; // @[LZD.scala 39:30]
  wire  _T_11; // @[LZD.scala 39:27]
  wire  _T_12; // @[LZD.scala 39:25]
  wire [1:0] _T_13; // @[Cat.scala 29:58]
  wire  _T_14; // @[LZD.scala 44:32]
  wire  _T_16; // @[Shift.scala 12:21]
  wire  _T_18; // @[LZD.scala 55:32]
  wire  _T_19; // @[LZD.scala 55:20]
  wire [1:0] _T_20; // @[Cat.scala 29:58]
  wire [1:0] _T_21; // @[convert.scala 21:22]
  wire [1:0] _T_22; // @[convert.scala 22:36]
  wire  _T_23; // @[Shift.scala 16:24]
  wire  _T_24; // @[Shift.scala 17:37]
  wire  _T_26; // @[Shift.scala 64:52]
  wire [1:0] _T_27; // @[Cat.scala 29:58]
  wire [1:0] _T_28; // @[Shift.scala 64:27]
  wire [1:0] _T_29; // @[Shift.scala 16:10]
  wire  _T_30; // @[convert.scala 23:34]
  wire  decA_fraction; // @[convert.scala 24:34]
  wire  _T_32; // @[convert.scala 25:26]
  wire [1:0] _T_34; // @[convert.scala 25:42]
  wire  _T_37; // @[convert.scala 26:67]
  wire  _T_38; // @[convert.scala 26:51]
  wire [3:0] _T_39; // @[Cat.scala 29:58]
  wire [3:0] _T_41; // @[convert.scala 29:56]
  wire  _T_42; // @[convert.scala 29:60]
  wire  _T_43; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_46; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [3:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_55; // @[convert.scala 18:24]
  wire  _T_56; // @[convert.scala 18:40]
  wire  _T_57; // @[convert.scala 18:36]
  wire [2:0] _T_58; // @[convert.scala 19:24]
  wire [2:0] _T_59; // @[convert.scala 19:43]
  wire [2:0] _T_60; // @[convert.scala 19:39]
  wire [1:0] _T_61; // @[LZD.scala 43:32]
  wire  _T_62; // @[LZD.scala 39:14]
  wire  _T_63; // @[LZD.scala 39:21]
  wire  _T_64; // @[LZD.scala 39:30]
  wire  _T_65; // @[LZD.scala 39:27]
  wire  _T_66; // @[LZD.scala 39:25]
  wire [1:0] _T_67; // @[Cat.scala 29:58]
  wire  _T_68; // @[LZD.scala 44:32]
  wire  _T_70; // @[Shift.scala 12:21]
  wire  _T_72; // @[LZD.scala 55:32]
  wire  _T_73; // @[LZD.scala 55:20]
  wire [1:0] _T_74; // @[Cat.scala 29:58]
  wire [1:0] _T_75; // @[convert.scala 21:22]
  wire [1:0] _T_76; // @[convert.scala 22:36]
  wire  _T_77; // @[Shift.scala 16:24]
  wire  _T_78; // @[Shift.scala 17:37]
  wire  _T_80; // @[Shift.scala 64:52]
  wire [1:0] _T_81; // @[Cat.scala 29:58]
  wire [1:0] _T_82; // @[Shift.scala 64:27]
  wire [1:0] _T_83; // @[Shift.scala 16:10]
  wire  _T_84; // @[convert.scala 23:34]
  wire  decB_fraction; // @[convert.scala 24:34]
  wire  _T_86; // @[convert.scala 25:26]
  wire [1:0] _T_88; // @[convert.scala 25:42]
  wire  _T_91; // @[convert.scala 26:67]
  wire  _T_92; // @[convert.scala 26:51]
  wire [3:0] _T_93; // @[Cat.scala 29:58]
  wire [3:0] _T_95; // @[convert.scala 29:56]
  wire  _T_96; // @[convert.scala 29:60]
  wire  _T_97; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_100; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [3:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_109; // @[Bitwise.scala 71:12]
  wire  _T_110; // @[PositDivisionSqrt.scala 80:40]
  wire [7:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_113; // @[PositDivisionSqrt.scala 82:31]
  wire [7:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_116; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_117; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_118; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_119; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_120; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_121; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_122; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_123; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_124; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_125; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [4:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_128; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_129; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_130; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_131; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_132; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_133; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_134; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_135; // @[PositDivisionSqrt.scala 117:30]
  wire [3:0] _T_137; // @[PositDivisionSqrt.scala 119:26]
  wire [3:0] _T_138; // @[PositDivisionSqrt.scala 118:20]
  wire [3:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [3:0] _T_139; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_141; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_142; // @[PositDivisionSqrt.scala 123:27]
  wire [2:0] _T_144; // @[PositDivisionSqrt.scala 123:52]
  wire [2:0] _T_145; // @[PositDivisionSqrt.scala 123:20]
  wire [3:0] _GEN_10; // @[PositDivisionSqrt.scala 122:64]
  wire [3:0] _T_146; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_148; // @[PositDivisionSqrt.scala 124:27]
  wire [3:0] _GEN_11; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _T_150; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _GEN_0; // @[PositDivisionSqrt.scala 116:29]
  wire [2:0] _T_151; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_153; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_154; // @[PositDivisionSqrt.scala 137:28]
  wire [7:0] _T_155; // @[PositDivisionSqrt.scala 146:22]
  wire [5:0] _T_156; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_157; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_158; // @[PositDivisionSqrt.scala 148:23]
  wire [7:0] _T_159; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_160; // @[PositDivisionSqrt.scala 149:23]
  wire [8:0] _T_161; // @[PositDivisionSqrt.scala 149:46]
  wire [7:0] _T_162; // @[PositDivisionSqrt.scala 149:56]
  wire [7:0] _T_163; // @[PositDivisionSqrt.scala 149:16]
  wire [7:0] _T_164; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_165; // @[PositDivisionSqrt.scala 150:17]
  wire [7:0] _T_166; // @[PositDivisionSqrt.scala 150:16]
  wire [7:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_168; // @[PositDivisionSqrt.scala 152:29]
  wire [7:0] _T_169; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_170; // @[PositDivisionSqrt.scala 153:29]
  wire [4:0] _T_171; // @[PositDivisionSqrt.scala 153:22]
  wire [7:0] _GEN_12; // @[PositDivisionSqrt.scala 152:93]
  wire [7:0] _T_172; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_174; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_175; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_176; // @[PositDivisionSqrt.scala 154:57]
  wire [7:0] _T_179; // @[Cat.scala 29:58]
  wire [7:0] _T_180; // @[PositDivisionSqrt.scala 154:22]
  wire [7:0] _T_181; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_183; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_184; // @[PositDivisionSqrt.scala 156:83]
  wire [3:0] _T_186; // @[Bitwise.scala 71:12]
  wire [6:0] bitMask; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  wire [6:0] _GEN_13; // @[PositDivisionSqrt.scala 156:53]
  wire [6:0] _T_187; // @[PositDivisionSqrt.scala 156:53]
  wire [7:0] _GEN_14; // @[PositDivisionSqrt.scala 155:51]
  wire [7:0] _T_188; // @[PositDivisionSqrt.scala 155:51]
  wire [5:0] _T_189; // @[PositDivisionSqrt.scala 157:53]
  wire [7:0] _GEN_15; // @[PositDivisionSqrt.scala 156:89]
  wire [7:0] _T_190; // @[PositDivisionSqrt.scala 156:89]
  wire [7:0] _T_191; // @[PositDivisionSqrt.scala 155:22]
  wire [7:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_193; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_194; // @[PositDivisionSqrt.scala 162:40]
  wire [7:0] _T_197; // @[PositDivisionSqrt.scala 163:97]
  wire [7:0] _T_199; // @[PositDivisionSqrt.scala 164:97]
  wire [7:0] _T_200; // @[PositDivisionSqrt.scala 161:92]
  wire [8:0] _T_205; // @[PositDivisionSqrt.scala 168:98]
  wire [7:0] _T_206; // @[PositDivisionSqrt.scala 168:108]
  wire [7:0] _T_208; // @[PositDivisionSqrt.scala 168:112]
  wire [7:0] _T_212; // @[PositDivisionSqrt.scala 169:112]
  wire [7:0] _T_213; // @[PositDivisionSqrt.scala 166:26]
  wire [7:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_214; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_215; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_217; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_218; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_219; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_220; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_221; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_223; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_224; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_225; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_226; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_227; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_230; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_231; // @[PositDivisionSqrt.scala 187:28]
  wire [7:0] _T_234; // @[PositDivisionSqrt.scala 188:47]
  wire [7:0] _T_235; // @[PositDivisionSqrt.scala 188:18]
  wire [5:0] _T_237; // @[PositDivisionSqrt.scala 189:18]
  wire [7:0] _GEN_16; // @[PositDivisionSqrt.scala 188:78]
  wire [7:0] _T_238; // @[PositDivisionSqrt.scala 188:78]
  wire [7:0] _GEN_17; // @[PositDivisionSqrt.scala 190:47]
  wire [7:0] _T_240; // @[PositDivisionSqrt.scala 190:47]
  wire [7:0] _T_241; // @[PositDivisionSqrt.scala 190:18]
  wire [7:0] _T_242; // @[PositDivisionSqrt.scala 189:78]
  wire [1:0] _T_244; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [7:0] _GEN_18; // @[PositDivisionSqrt.scala 197:25]
  wire [7:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire  _T_247; // @[PositDivisionSqrt.scala 200:97]
  wire  _T_248; // @[PositDivisionSqrt.scala 201:97]
  wire  realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_249; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_250; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_251; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_254; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_255; // @[Cat.scala 29:58]
  wire [2:0] _T_256; // @[PositDivisionSqrt.scala 209:63]
  wire [4:0] _GEN_19; // @[PositDivisionSqrt.scala 209:31]
  wire [4:0] _T_258; // @[PositDivisionSqrt.scala 209:31]
  wire [4:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [4:0] _T_260; // @[Mux.scala 87:16]
  wire [4:0] _T_261; // @[Mux.scala 87:16]
  wire [2:0] _T_262; // @[PositDivisionSqrt.scala 224:48]
  wire [2:0] _T_263; // @[PositDivisionSqrt.scala 224:64]
  wire [2:0] decQ_grs; // @[PositDivisionSqrt.scala 224:23]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [3:0] _GEN_20; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [3:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire  _T_269; // @[convert.scala 46:61]
  wire  _T_270; // @[convert.scala 46:52]
  wire  _T_272; // @[convert.scala 46:42]
  wire [2:0] _T_273; // @[convert.scala 48:34]
  wire  _T_274; // @[convert.scala 49:36]
  wire [2:0] _T_276; // @[convert.scala 50:36]
  wire [2:0] _T_277; // @[convert.scala 50:36]
  wire [2:0] _T_278; // @[convert.scala 50:28]
  wire  _T_279; // @[convert.scala 51:31]
  wire  _T_280; // @[convert.scala 52:43]
  wire [6:0] _T_284; // @[Cat.scala 29:58]
  wire [2:0] _T_285; // @[Shift.scala 39:17]
  wire  _T_286; // @[Shift.scala 39:24]
  wire [2:0] _T_288; // @[Shift.scala 90:30]
  wire [3:0] _T_289; // @[Shift.scala 90:48]
  wire  _T_290; // @[Shift.scala 90:57]
  wire [2:0] _GEN_21; // @[Shift.scala 90:39]
  wire [2:0] _T_291; // @[Shift.scala 90:39]
  wire  _T_292; // @[Shift.scala 12:21]
  wire  _T_293; // @[Shift.scala 12:21]
  wire [3:0] _T_295; // @[Bitwise.scala 71:12]
  wire [6:0] _T_296; // @[Cat.scala 29:58]
  wire [6:0] _T_297; // @[Shift.scala 91:22]
  wire [1:0] _T_298; // @[Shift.scala 92:77]
  wire [4:0] _T_299; // @[Shift.scala 90:30]
  wire [1:0] _T_300; // @[Shift.scala 90:48]
  wire  _T_301; // @[Shift.scala 90:57]
  wire [4:0] _GEN_22; // @[Shift.scala 90:39]
  wire [4:0] _T_302; // @[Shift.scala 90:39]
  wire  _T_303; // @[Shift.scala 12:21]
  wire  _T_304; // @[Shift.scala 12:21]
  wire [1:0] _T_306; // @[Bitwise.scala 71:12]
  wire [6:0] _T_307; // @[Cat.scala 29:58]
  wire [6:0] _T_308; // @[Shift.scala 91:22]
  wire  _T_309; // @[Shift.scala 92:77]
  wire [5:0] _T_310; // @[Shift.scala 90:30]
  wire  _T_311; // @[Shift.scala 90:48]
  wire [5:0] _GEN_23; // @[Shift.scala 90:39]
  wire [5:0] _T_313; // @[Shift.scala 90:39]
  wire  _T_315; // @[Shift.scala 12:21]
  wire [6:0] _T_316; // @[Cat.scala 29:58]
  wire [6:0] _T_317; // @[Shift.scala 91:22]
  wire [6:0] _T_320; // @[Bitwise.scala 71:12]
  wire [6:0] _T_321; // @[Shift.scala 39:10]
  wire  _T_322; // @[convert.scala 55:31]
  wire  _T_323; // @[convert.scala 56:31]
  wire  _T_324; // @[convert.scala 57:31]
  wire  _T_325; // @[convert.scala 58:31]
  wire [3:0] _T_326; // @[convert.scala 59:69]
  wire  _T_327; // @[convert.scala 59:81]
  wire  _T_328; // @[convert.scala 59:50]
  wire  _T_330; // @[convert.scala 60:81]
  wire  _T_331; // @[convert.scala 61:44]
  wire  _T_332; // @[convert.scala 61:52]
  wire  _T_333; // @[convert.scala 61:36]
  wire  _T_334; // @[convert.scala 62:63]
  wire  _T_335; // @[convert.scala 62:103]
  wire  _T_336; // @[convert.scala 62:60]
  wire [3:0] _GEN_24; // @[convert.scala 63:56]
  wire [3:0] _T_339; // @[convert.scala 63:56]
  wire [4:0] _T_340; // @[Cat.scala 29:58]
  wire [4:0] _T_342; // @[Mux.scala 87:16]
  assign _T_1 = io_A[4]; // @[convert.scala 18:24]
  assign _T_2 = io_A[3]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[3:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[2:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[2:1]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7 != 2'h0; // @[LZD.scala 39:14]
  assign _T_9 = _T_7[1]; // @[LZD.scala 39:21]
  assign _T_10 = _T_7[0]; // @[LZD.scala 39:30]
  assign _T_11 = ~ _T_10; // @[LZD.scala 39:27]
  assign _T_12 = _T_9 | _T_11; // @[LZD.scala 39:25]
  assign _T_13 = {_T_8,_T_12}; // @[Cat.scala 29:58]
  assign _T_14 = _T_6[0:0]; // @[LZD.scala 44:32]
  assign _T_16 = _T_13[1]; // @[Shift.scala 12:21]
  assign _T_18 = _T_13[0:0]; // @[LZD.scala 55:32]
  assign _T_19 = _T_16 ? _T_18 : _T_14; // @[LZD.scala 55:20]
  assign _T_20 = {_T_16,_T_19}; // @[Cat.scala 29:58]
  assign _T_21 = ~ _T_20; // @[convert.scala 21:22]
  assign _T_22 = io_A[1:0]; // @[convert.scala 22:36]
  assign _T_23 = _T_21 < 2'h2; // @[Shift.scala 16:24]
  assign _T_24 = _T_21[0]; // @[Shift.scala 17:37]
  assign _T_26 = _T_22[0:0]; // @[Shift.scala 64:52]
  assign _T_27 = {_T_26,1'h0}; // @[Cat.scala 29:58]
  assign _T_28 = _T_24 ? _T_27 : _T_22; // @[Shift.scala 64:27]
  assign _T_29 = _T_23 ? _T_28 : 2'h0; // @[Shift.scala 16:10]
  assign _T_30 = _T_29[1:1]; // @[convert.scala 23:34]
  assign decA_fraction = _T_29[0:0]; // @[convert.scala 24:34]
  assign _T_32 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_34 = _T_3 ? _T_21 : _T_20; // @[convert.scala 25:42]
  assign _T_37 = ~ _T_30; // @[convert.scala 26:67]
  assign _T_38 = _T_1 ? _T_37 : _T_30; // @[convert.scala 26:51]
  assign _T_39 = {_T_32,_T_34,_T_38}; // @[Cat.scala 29:58]
  assign _T_41 = io_A[3:0]; // @[convert.scala 29:56]
  assign _T_42 = _T_41 != 4'h0; // @[convert.scala 29:60]
  assign _T_43 = ~ _T_42; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_43; // @[convert.scala 29:39]
  assign _T_46 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_46 & _T_43; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_39); // @[convert.scala 32:24]
  assign _T_55 = io_B[4]; // @[convert.scala 18:24]
  assign _T_56 = io_B[3]; // @[convert.scala 18:40]
  assign _T_57 = _T_55 ^ _T_56; // @[convert.scala 18:36]
  assign _T_58 = io_B[3:1]; // @[convert.scala 19:24]
  assign _T_59 = io_B[2:0]; // @[convert.scala 19:43]
  assign _T_60 = _T_58 ^ _T_59; // @[convert.scala 19:39]
  assign _T_61 = _T_60[2:1]; // @[LZD.scala 43:32]
  assign _T_62 = _T_61 != 2'h0; // @[LZD.scala 39:14]
  assign _T_63 = _T_61[1]; // @[LZD.scala 39:21]
  assign _T_64 = _T_61[0]; // @[LZD.scala 39:30]
  assign _T_65 = ~ _T_64; // @[LZD.scala 39:27]
  assign _T_66 = _T_63 | _T_65; // @[LZD.scala 39:25]
  assign _T_67 = {_T_62,_T_66}; // @[Cat.scala 29:58]
  assign _T_68 = _T_60[0:0]; // @[LZD.scala 44:32]
  assign _T_70 = _T_67[1]; // @[Shift.scala 12:21]
  assign _T_72 = _T_67[0:0]; // @[LZD.scala 55:32]
  assign _T_73 = _T_70 ? _T_72 : _T_68; // @[LZD.scala 55:20]
  assign _T_74 = {_T_70,_T_73}; // @[Cat.scala 29:58]
  assign _T_75 = ~ _T_74; // @[convert.scala 21:22]
  assign _T_76 = io_B[1:0]; // @[convert.scala 22:36]
  assign _T_77 = _T_75 < 2'h2; // @[Shift.scala 16:24]
  assign _T_78 = _T_75[0]; // @[Shift.scala 17:37]
  assign _T_80 = _T_76[0:0]; // @[Shift.scala 64:52]
  assign _T_81 = {_T_80,1'h0}; // @[Cat.scala 29:58]
  assign _T_82 = _T_78 ? _T_81 : _T_76; // @[Shift.scala 64:27]
  assign _T_83 = _T_77 ? _T_82 : 2'h0; // @[Shift.scala 16:10]
  assign _T_84 = _T_83[1:1]; // @[convert.scala 23:34]
  assign decB_fraction = _T_83[0:0]; // @[convert.scala 24:34]
  assign _T_86 = _T_57 == 1'h0; // @[convert.scala 25:26]
  assign _T_88 = _T_57 ? _T_75 : _T_74; // @[convert.scala 25:42]
  assign _T_91 = ~ _T_84; // @[convert.scala 26:67]
  assign _T_92 = _T_55 ? _T_91 : _T_84; // @[convert.scala 26:51]
  assign _T_93 = {_T_86,_T_88,_T_92}; // @[Cat.scala 29:58]
  assign _T_95 = io_B[3:0]; // @[convert.scala 29:56]
  assign _T_96 = _T_95 != 4'h0; // @[convert.scala 29:60]
  assign _T_97 = ~ _T_96; // @[convert.scala 29:41]
  assign decB_isNaR = _T_55 & _T_97; // @[convert.scala 29:39]
  assign _T_100 = _T_55 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_100 & _T_97; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_93); // @[convert.scala 32:24]
  assign _T_109 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_110 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_109,_T_110,decA_fraction,3'h0}; // @[Cat.scala 29:58]
  assign _T_113 = ~ _T_55; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_55,_T_113,decB_fraction,5'h0}; // @[Cat.scala 29:58]
  assign _T_116 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_116 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_117 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_118 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_119 = _T_118 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_120 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_121 = decA_isZero & _T_120; // @[PositDivisionSqrt.scala 94:43]
  assign _T_122 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_123 = _T_121 & _T_122; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_124 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_125 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_124 & _T_125; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_124 & _T_46; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_128 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_128; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 3'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 3'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_129 = sigX_Z[7]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_130 = sigX_Z[5]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_129 ^ _T_130; // @[PositDivisionSqrt.scala 113:50]
  assign _T_131 = cycleNum == 3'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_131 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_132 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_133 = _T_132 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_134 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_135 = entering & _T_134; // @[PositDivisionSqrt.scala 117:30]
  assign _T_137 = io_sqrtOp ? 4'h6 : 4'h8; // @[PositDivisionSqrt.scala 119:26]
  assign _T_138 = entering_normalCase ? _T_137 : 4'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{3'd0}, _T_135}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_139 = _GEN_9 | _T_138; // @[PositDivisionSqrt.scala 117:64]
  assign _T_141 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_142 = _T_132 & _T_141; // @[PositDivisionSqrt.scala 123:27]
  assign _T_144 = cycleNum - 3'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_145 = _T_142 ? _T_144 : 3'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _GEN_10 = {{1'd0}, _T_145}; // @[PositDivisionSqrt.scala 122:64]
  assign _T_146 = _T_139 | _GEN_10; // @[PositDivisionSqrt.scala 122:64]
  assign _T_148 = _T_132 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_11 = {{3'd0}, _T_148}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_150 = _T_146 | _GEN_11; // @[PositDivisionSqrt.scala 123:64]
  assign _GEN_0 = _T_133 ? _T_150 : {{1'd0}, cycleNum}; // @[PositDivisionSqrt.scala 116:29]
  assign _T_151 = decA_scale[3:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_153 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_154 = entering_normalCase & _T_153; // @[PositDivisionSqrt.scala 137:28]
  assign _T_155 = 8'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign _T_156 = _T_155[7:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_157 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_158 = ready & _T_157; // @[PositDivisionSqrt.scala 148:23]
  assign _T_159 = _T_158 ? sigA_S : 8'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_160 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_161 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_162 = _T_161[7:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_163 = _T_160 ? _T_162 : 8'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_164 = _T_159 | _T_163; // @[PositDivisionSqrt.scala 148:66]
  assign _T_165 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_166 = _T_165 ? rem_Z : 8'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_164 | _T_166; // @[PositDivisionSqrt.scala 149:66]
  assign _T_168 = ready & _T_153; // @[PositDivisionSqrt.scala 152:29]
  assign _T_169 = _T_168 ? sigB_S : 8'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_170 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_171 = _T_170 ? 5'h10 : 5'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_12 = {{3'd0}, _T_171}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_172 = _T_169 | _GEN_12; // @[PositDivisionSqrt.scala 152:93]
  assign _T_174 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_175 = _T_165 & _T_174; // @[PositDivisionSqrt.scala 154:30]
  assign _T_176 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_179 = {signB_Z,_T_176,fractB_Z,5'h0}; // @[Cat.scala 29:58]
  assign _T_180 = _T_175 ? _T_179 : 8'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_181 = _T_172 | _T_180; // @[PositDivisionSqrt.scala 153:93]
  assign _T_183 = _T_165 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_184 = rem[7:7]; // @[PositDivisionSqrt.scala 156:83]
  assign _T_186 = _T_184 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign bitMask = {{1'd0}, _T_156}; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  assign _GEN_13 = {{3'd0}, _T_186}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_187 = bitMask & _GEN_13; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_14 = {{1'd0}, _T_187}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_188 = sigX_Z | _GEN_14; // @[PositDivisionSqrt.scala 155:51]
  assign _T_189 = bitMask[6:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_15 = {{2'd0}, _T_189}; // @[PositDivisionSqrt.scala 156:89]
  assign _T_190 = _T_188 | _GEN_15; // @[PositDivisionSqrt.scala 156:89]
  assign _T_191 = _T_183 ? _T_190 : 8'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_181 | _T_191; // @[PositDivisionSqrt.scala 154:93]
  assign _T_193 = trialTerm[7:7]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_194 = _T_184 ^ _T_193; // @[PositDivisionSqrt.scala 162:40]
  assign _T_197 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_199 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_200 = _T_194 ? _T_197 : _T_199; // @[PositDivisionSqrt.scala 161:92]
  assign _T_205 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_206 = _T_205[7:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_208 = _T_206 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_212 = _T_206 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_213 = _T_194 ? _T_208 : _T_212; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_200 : _T_213; // @[PositDivisionSqrt.scala 159:27]
  assign _T_214 = trialRem != 8'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_214 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_215 = rem != 8'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_215 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_217 = trialRem[7:7]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_218 = _T_193 ^ _T_217; // @[PositDivisionSqrt.scala 176:49]
  assign _T_219 = ~ _T_218; // @[PositDivisionSqrt.scala 176:29]
  assign _T_220 = sigX_Z[7:7]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_221 = ~ _T_220; // @[PositDivisionSqrt.scala 178:49]
  assign _T_223 = remIsZero ? _T_220 : _T_219; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_221 : _T_223; // @[Mux.scala 87:16]
  assign _T_224 = cycleNum > 3'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_225 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_226 = _T_224 & _T_225; // @[PositDivisionSqrt.scala 183:48]
  assign _T_227 = entering_normalCase | _T_226; // @[PositDivisionSqrt.scala 183:28]
  assign _T_230 = _T_165 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_231 = entering_normalCase | _T_230; // @[PositDivisionSqrt.scala 187:28]
  assign _T_234 = {newBit, 7'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_235 = _T_168 ? _T_234 : 8'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_237 = _T_170 ? 6'h20 : 6'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_16 = {{2'd0}, _T_237}; // @[PositDivisionSqrt.scala 188:78]
  assign _T_238 = _T_235 | _GEN_16; // @[PositDivisionSqrt.scala 188:78]
  assign _GEN_17 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_240 = sigX_Z | _GEN_17; // @[PositDivisionSqrt.scala 190:47]
  assign _T_241 = _T_165 ? _T_240 : 8'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_242 = _T_238 | _T_241; // @[PositDivisionSqrt.scala 189:78]
  assign _T_244 = {_T_220, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_244 : {{1'd0}, _T_220}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_18 = {{6'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_18; // @[PositDivisionSqrt.scala 197:25]
  assign _T_247 = realSigX[4]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_248 = realSigX[3]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_247 : _T_248; // @[PositDivisionSqrt.scala 198:21]
  assign _T_249 = realSigX[7]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_250 = realSigX[5]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_251 = _T_249 ^ _T_250; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_251; // @[PositDivisionSqrt.scala 205:23]
  assign notNeedSubTwo = _T_249 ^ _T_247; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_254 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_254; // @[PositDivisionSqrt.scala 208:36]
  assign _T_255 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_256 = {1'b0,$signed(_T_255)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_19 = {{2{_T_256[2]}},_T_256}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_258 = $signed(scale_Z) - $signed(_GEN_19); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_258); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-5'sh7); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(5'sh6); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[7:7]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_260 = underflow ? $signed(-5'sh7) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_261 = overflow ? $signed(5'sh6) : $signed(_T_260); // @[Mux.scala 87:16]
  assign _T_262 = realSigX[3:1]; // @[PositDivisionSqrt.scala 224:48]
  assign _T_263 = realSigX[2:0]; // @[PositDivisionSqrt.scala 224:64]
  assign decQ_grs = scaleNotChange ? _T_262 : _T_263; // @[PositDivisionSqrt.scala 224:23]
  assign outValid = cycleNum == 3'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_20 = _T_261[3:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_20); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_269 = decQ_scale[0]; // @[convert.scala 46:61]
  assign _T_270 = ~ _T_269; // @[convert.scala 46:52]
  assign _T_272 = decQ_sign ? _T_270 : _T_269; // @[convert.scala 46:42]
  assign _T_273 = decQ_scale[3:1]; // @[convert.scala 48:34]
  assign _T_274 = _T_273[2:2]; // @[convert.scala 49:36]
  assign _T_276 = ~ _T_273; // @[convert.scala 50:36]
  assign _T_277 = $signed(_T_276); // @[convert.scala 50:36]
  assign _T_278 = _T_274 ? $signed(_T_277) : $signed(_T_273); // @[convert.scala 50:28]
  assign _T_279 = _T_274 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_280 = ~ _T_279; // @[convert.scala 52:43]
  assign _T_284 = {_T_280,_T_279,_T_272,realFrac,decQ_grs}; // @[Cat.scala 29:58]
  assign _T_285 = $unsigned(_T_278); // @[Shift.scala 39:17]
  assign _T_286 = _T_285 < 3'h7; // @[Shift.scala 39:24]
  assign _T_288 = _T_284[6:4]; // @[Shift.scala 90:30]
  assign _T_289 = _T_284[3:0]; // @[Shift.scala 90:48]
  assign _T_290 = _T_289 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{2'd0}, _T_290}; // @[Shift.scala 90:39]
  assign _T_291 = _T_288 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_292 = _T_285[2]; // @[Shift.scala 12:21]
  assign _T_293 = _T_284[6]; // @[Shift.scala 12:21]
  assign _T_295 = _T_293 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_296 = {_T_295,_T_291}; // @[Cat.scala 29:58]
  assign _T_297 = _T_292 ? _T_296 : _T_284; // @[Shift.scala 91:22]
  assign _T_298 = _T_285[1:0]; // @[Shift.scala 92:77]
  assign _T_299 = _T_297[6:2]; // @[Shift.scala 90:30]
  assign _T_300 = _T_297[1:0]; // @[Shift.scala 90:48]
  assign _T_301 = _T_300 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{4'd0}, _T_301}; // @[Shift.scala 90:39]
  assign _T_302 = _T_299 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_303 = _T_298[1]; // @[Shift.scala 12:21]
  assign _T_304 = _T_297[6]; // @[Shift.scala 12:21]
  assign _T_306 = _T_304 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_307 = {_T_306,_T_302}; // @[Cat.scala 29:58]
  assign _T_308 = _T_303 ? _T_307 : _T_297; // @[Shift.scala 91:22]
  assign _T_309 = _T_298[0:0]; // @[Shift.scala 92:77]
  assign _T_310 = _T_308[6:1]; // @[Shift.scala 90:30]
  assign _T_311 = _T_308[0:0]; // @[Shift.scala 90:48]
  assign _GEN_23 = {{5'd0}, _T_311}; // @[Shift.scala 90:39]
  assign _T_313 = _T_310 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_315 = _T_308[6]; // @[Shift.scala 12:21]
  assign _T_316 = {_T_315,_T_313}; // @[Cat.scala 29:58]
  assign _T_317 = _T_309 ? _T_316 : _T_308; // @[Shift.scala 91:22]
  assign _T_320 = _T_293 ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign _T_321 = _T_286 ? _T_317 : _T_320; // @[Shift.scala 39:10]
  assign _T_322 = _T_321[3]; // @[convert.scala 55:31]
  assign _T_323 = _T_321[2]; // @[convert.scala 56:31]
  assign _T_324 = _T_321[1]; // @[convert.scala 57:31]
  assign _T_325 = _T_321[0]; // @[convert.scala 58:31]
  assign _T_326 = _T_321[6:3]; // @[convert.scala 59:69]
  assign _T_327 = _T_326 != 4'h0; // @[convert.scala 59:81]
  assign _T_328 = ~ _T_327; // @[convert.scala 59:50]
  assign _T_330 = _T_326 == 4'hf; // @[convert.scala 60:81]
  assign _T_331 = _T_322 | _T_324; // @[convert.scala 61:44]
  assign _T_332 = _T_331 | _T_325; // @[convert.scala 61:52]
  assign _T_333 = _T_323 & _T_332; // @[convert.scala 61:36]
  assign _T_334 = ~ _T_330; // @[convert.scala 62:63]
  assign _T_335 = _T_334 & _T_333; // @[convert.scala 62:103]
  assign _T_336 = _T_328 | _T_335; // @[convert.scala 62:60]
  assign _GEN_24 = {{3'd0}, _T_336}; // @[convert.scala 63:56]
  assign _T_339 = _T_326 + _GEN_24; // @[convert.scala 63:56]
  assign _T_340 = {decQ_sign,_T_339}; // @[Cat.scala 29:58]
  assign _T_342 = isZero_Z ? 5'h0 : _T_340; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 3'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_174; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 5'h10 : _T_342; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 3'h0;
    end else begin
      cycleNum <= _GEN_0[2:0];
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_117;
      end else begin
        isNaR_Z <= _T_119;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_123;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_151[2]}},_T_151};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_154) begin
      signB_Z <= _T_55;
    end
    if (_T_154) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_227) begin
      if (ready) begin
        if (_T_194) begin
          rem_Z <= _T_197;
        end else begin
          rem_Z <= _T_199;
        end
      end else begin
        if (_T_194) begin
          rem_Z <= _T_208;
        end else begin
          rem_Z <= _T_212;
        end
      end
    end
    if (_T_231) begin
      sigX_Z <= _T_242;
    end
  end
endmodule
