module FMA_Dec5_1(
  input        clock,
  input        reset,
  input  [4:0] io_A,
  input  [4:0] io_B,
  input  [4:0] io_C,
  output [2:0] io_sigA,
  output [2:0] io_sigB,
  output       io_outIsNaR,
  output       io_Csign,
  output       io_CisNar,
  output       io_CisZero,
  output       io_Cfrac,
  output [3:0] io_Ascale,
  output [3:0] io_Bscale,
  output [3:0] io_Cscale
);
  wire [5:0] _T_2; // @[FMA_Dec.scala 38:46]
  wire [4:0] realA; // @[FMA_Dec.scala 38:46]
  wire [5:0] _T_5; // @[FMA_Dec.scala 39:46]
  wire [4:0] realC; // @[FMA_Dec.scala 39:46]
  wire  _T_7; // @[convert.scala 18:24]
  wire  _T_8; // @[convert.scala 18:40]
  wire  _T_9; // @[convert.scala 18:36]
  wire [2:0] _T_10; // @[convert.scala 19:24]
  wire [2:0] _T_11; // @[convert.scala 19:43]
  wire [2:0] _T_12; // @[convert.scala 19:39]
  wire [1:0] _T_13; // @[LZD.scala 43:32]
  wire  _T_14; // @[LZD.scala 39:14]
  wire  _T_15; // @[LZD.scala 39:21]
  wire  _T_16; // @[LZD.scala 39:30]
  wire  _T_17; // @[LZD.scala 39:27]
  wire  _T_18; // @[LZD.scala 39:25]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  _T_20; // @[LZD.scala 44:32]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_24; // @[LZD.scala 55:32]
  wire  _T_25; // @[LZD.scala 55:20]
  wire [1:0] _T_26; // @[Cat.scala 29:58]
  wire [1:0] _T_27; // @[convert.scala 21:22]
  wire [1:0] _T_28; // @[convert.scala 22:36]
  wire  _T_29; // @[Shift.scala 16:24]
  wire  _T_30; // @[Shift.scala 17:37]
  wire  _T_32; // @[Shift.scala 64:52]
  wire [1:0] _T_33; // @[Cat.scala 29:58]
  wire [1:0] _T_34; // @[Shift.scala 64:27]
  wire [1:0] _T_35; // @[Shift.scala 16:10]
  wire  _T_36; // @[convert.scala 23:34]
  wire  decA_fraction; // @[convert.scala 24:34]
  wire  _T_38; // @[convert.scala 25:26]
  wire [1:0] _T_40; // @[convert.scala 25:42]
  wire  _T_43; // @[convert.scala 26:67]
  wire  _T_44; // @[convert.scala 26:51]
  wire [3:0] _T_45; // @[Cat.scala 29:58]
  wire [3:0] _T_47; // @[convert.scala 29:56]
  wire  _T_48; // @[convert.scala 29:60]
  wire  _T_49; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_52; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire  _T_61; // @[convert.scala 18:24]
  wire  _T_62; // @[convert.scala 18:40]
  wire  _T_63; // @[convert.scala 18:36]
  wire [2:0] _T_64; // @[convert.scala 19:24]
  wire [2:0] _T_65; // @[convert.scala 19:43]
  wire [2:0] _T_66; // @[convert.scala 19:39]
  wire [1:0] _T_67; // @[LZD.scala 43:32]
  wire  _T_68; // @[LZD.scala 39:14]
  wire  _T_69; // @[LZD.scala 39:21]
  wire  _T_70; // @[LZD.scala 39:30]
  wire  _T_71; // @[LZD.scala 39:27]
  wire  _T_72; // @[LZD.scala 39:25]
  wire [1:0] _T_73; // @[Cat.scala 29:58]
  wire  _T_74; // @[LZD.scala 44:32]
  wire  _T_76; // @[Shift.scala 12:21]
  wire  _T_78; // @[LZD.scala 55:32]
  wire  _T_79; // @[LZD.scala 55:20]
  wire [1:0] _T_80; // @[Cat.scala 29:58]
  wire [1:0] _T_81; // @[convert.scala 21:22]
  wire [1:0] _T_82; // @[convert.scala 22:36]
  wire  _T_83; // @[Shift.scala 16:24]
  wire  _T_84; // @[Shift.scala 17:37]
  wire  _T_86; // @[Shift.scala 64:52]
  wire [1:0] _T_87; // @[Cat.scala 29:58]
  wire [1:0] _T_88; // @[Shift.scala 64:27]
  wire [1:0] _T_89; // @[Shift.scala 16:10]
  wire  _T_90; // @[convert.scala 23:34]
  wire  decB_fraction; // @[convert.scala 24:34]
  wire  _T_92; // @[convert.scala 25:26]
  wire [1:0] _T_94; // @[convert.scala 25:42]
  wire  _T_97; // @[convert.scala 26:67]
  wire  _T_98; // @[convert.scala 26:51]
  wire [3:0] _T_99; // @[Cat.scala 29:58]
  wire [3:0] _T_101; // @[convert.scala 29:56]
  wire  _T_102; // @[convert.scala 29:60]
  wire  _T_103; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_106; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire  _T_115; // @[convert.scala 18:24]
  wire  _T_116; // @[convert.scala 18:40]
  wire  _T_117; // @[convert.scala 18:36]
  wire [2:0] _T_118; // @[convert.scala 19:24]
  wire [2:0] _T_119; // @[convert.scala 19:43]
  wire [2:0] _T_120; // @[convert.scala 19:39]
  wire [1:0] _T_121; // @[LZD.scala 43:32]
  wire  _T_122; // @[LZD.scala 39:14]
  wire  _T_123; // @[LZD.scala 39:21]
  wire  _T_124; // @[LZD.scala 39:30]
  wire  _T_125; // @[LZD.scala 39:27]
  wire  _T_126; // @[LZD.scala 39:25]
  wire [1:0] _T_127; // @[Cat.scala 29:58]
  wire  _T_128; // @[LZD.scala 44:32]
  wire  _T_130; // @[Shift.scala 12:21]
  wire  _T_132; // @[LZD.scala 55:32]
  wire  _T_133; // @[LZD.scala 55:20]
  wire [1:0] _T_134; // @[Cat.scala 29:58]
  wire [1:0] _T_135; // @[convert.scala 21:22]
  wire [1:0] _T_136; // @[convert.scala 22:36]
  wire  _T_137; // @[Shift.scala 16:24]
  wire  _T_138; // @[Shift.scala 17:37]
  wire  _T_140; // @[Shift.scala 64:52]
  wire [1:0] _T_141; // @[Cat.scala 29:58]
  wire [1:0] _T_142; // @[Shift.scala 64:27]
  wire [1:0] _T_143; // @[Shift.scala 16:10]
  wire  _T_144; // @[convert.scala 23:34]
  wire  _T_146; // @[convert.scala 25:26]
  wire [1:0] _T_148; // @[convert.scala 25:42]
  wire  _T_151; // @[convert.scala 26:67]
  wire  _T_152; // @[convert.scala 26:51]
  wire [3:0] _T_153; // @[Cat.scala 29:58]
  wire [3:0] _T_155; // @[convert.scala 29:56]
  wire  _T_156; // @[convert.scala 29:60]
  wire  _T_157; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_160; // @[convert.scala 30:19]
  wire  _T_168; // @[FMA_Dec.scala 46:30]
  wire  _T_170; // @[FMA_Dec.scala 49:34]
  wire  _T_171; // @[FMA_Dec.scala 49:47]
  wire  _T_172; // @[FMA_Dec.scala 49:45]
  wire [2:0] _T_174; // @[Cat.scala 29:58]
  wire  _T_176; // @[FMA_Dec.scala 50:34]
  wire  _T_177; // @[FMA_Dec.scala 50:47]
  wire  _T_178; // @[FMA_Dec.scala 50:45]
  wire [2:0] _T_180; // @[Cat.scala 29:58]
  assign _T_2 = {{1'd0}, io_A}; // @[FMA_Dec.scala 38:46]
  assign realA = _T_2[4:0]; // @[FMA_Dec.scala 38:46]
  assign _T_5 = {{1'd0}, io_C}; // @[FMA_Dec.scala 39:46]
  assign realC = _T_5[4:0]; // @[FMA_Dec.scala 39:46]
  assign _T_7 = realA[4]; // @[convert.scala 18:24]
  assign _T_8 = realA[3]; // @[convert.scala 18:40]
  assign _T_9 = _T_7 ^ _T_8; // @[convert.scala 18:36]
  assign _T_10 = realA[3:1]; // @[convert.scala 19:24]
  assign _T_11 = realA[2:0]; // @[convert.scala 19:43]
  assign _T_12 = _T_10 ^ _T_11; // @[convert.scala 19:39]
  assign _T_13 = _T_12[2:1]; // @[LZD.scala 43:32]
  assign _T_14 = _T_13 != 2'h0; // @[LZD.scala 39:14]
  assign _T_15 = _T_13[1]; // @[LZD.scala 39:21]
  assign _T_16 = _T_13[0]; // @[LZD.scala 39:30]
  assign _T_17 = ~ _T_16; // @[LZD.scala 39:27]
  assign _T_18 = _T_15 | _T_17; // @[LZD.scala 39:25]
  assign _T_19 = {_T_14,_T_18}; // @[Cat.scala 29:58]
  assign _T_20 = _T_12[0:0]; // @[LZD.scala 44:32]
  assign _T_22 = _T_19[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_19[0:0]; // @[LZD.scala 55:32]
  assign _T_25 = _T_22 ? _T_24 : _T_20; // @[LZD.scala 55:20]
  assign _T_26 = {_T_22,_T_25}; // @[Cat.scala 29:58]
  assign _T_27 = ~ _T_26; // @[convert.scala 21:22]
  assign _T_28 = realA[1:0]; // @[convert.scala 22:36]
  assign _T_29 = _T_27 < 2'h2; // @[Shift.scala 16:24]
  assign _T_30 = _T_27[0]; // @[Shift.scala 17:37]
  assign _T_32 = _T_28[0:0]; // @[Shift.scala 64:52]
  assign _T_33 = {_T_32,1'h0}; // @[Cat.scala 29:58]
  assign _T_34 = _T_30 ? _T_33 : _T_28; // @[Shift.scala 64:27]
  assign _T_35 = _T_29 ? _T_34 : 2'h0; // @[Shift.scala 16:10]
  assign _T_36 = _T_35[1:1]; // @[convert.scala 23:34]
  assign decA_fraction = _T_35[0:0]; // @[convert.scala 24:34]
  assign _T_38 = _T_9 == 1'h0; // @[convert.scala 25:26]
  assign _T_40 = _T_9 ? _T_27 : _T_26; // @[convert.scala 25:42]
  assign _T_43 = ~ _T_36; // @[convert.scala 26:67]
  assign _T_44 = _T_7 ? _T_43 : _T_36; // @[convert.scala 26:51]
  assign _T_45 = {_T_38,_T_40,_T_44}; // @[Cat.scala 29:58]
  assign _T_47 = realA[3:0]; // @[convert.scala 29:56]
  assign _T_48 = _T_47 != 4'h0; // @[convert.scala 29:60]
  assign _T_49 = ~ _T_48; // @[convert.scala 29:41]
  assign decA_isNaR = _T_7 & _T_49; // @[convert.scala 29:39]
  assign _T_52 = _T_7 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_52 & _T_49; // @[convert.scala 30:41]
  assign _T_61 = io_B[4]; // @[convert.scala 18:24]
  assign _T_62 = io_B[3]; // @[convert.scala 18:40]
  assign _T_63 = _T_61 ^ _T_62; // @[convert.scala 18:36]
  assign _T_64 = io_B[3:1]; // @[convert.scala 19:24]
  assign _T_65 = io_B[2:0]; // @[convert.scala 19:43]
  assign _T_66 = _T_64 ^ _T_65; // @[convert.scala 19:39]
  assign _T_67 = _T_66[2:1]; // @[LZD.scala 43:32]
  assign _T_68 = _T_67 != 2'h0; // @[LZD.scala 39:14]
  assign _T_69 = _T_67[1]; // @[LZD.scala 39:21]
  assign _T_70 = _T_67[0]; // @[LZD.scala 39:30]
  assign _T_71 = ~ _T_70; // @[LZD.scala 39:27]
  assign _T_72 = _T_69 | _T_71; // @[LZD.scala 39:25]
  assign _T_73 = {_T_68,_T_72}; // @[Cat.scala 29:58]
  assign _T_74 = _T_66[0:0]; // @[LZD.scala 44:32]
  assign _T_76 = _T_73[1]; // @[Shift.scala 12:21]
  assign _T_78 = _T_73[0:0]; // @[LZD.scala 55:32]
  assign _T_79 = _T_76 ? _T_78 : _T_74; // @[LZD.scala 55:20]
  assign _T_80 = {_T_76,_T_79}; // @[Cat.scala 29:58]
  assign _T_81 = ~ _T_80; // @[convert.scala 21:22]
  assign _T_82 = io_B[1:0]; // @[convert.scala 22:36]
  assign _T_83 = _T_81 < 2'h2; // @[Shift.scala 16:24]
  assign _T_84 = _T_81[0]; // @[Shift.scala 17:37]
  assign _T_86 = _T_82[0:0]; // @[Shift.scala 64:52]
  assign _T_87 = {_T_86,1'h0}; // @[Cat.scala 29:58]
  assign _T_88 = _T_84 ? _T_87 : _T_82; // @[Shift.scala 64:27]
  assign _T_89 = _T_83 ? _T_88 : 2'h0; // @[Shift.scala 16:10]
  assign _T_90 = _T_89[1:1]; // @[convert.scala 23:34]
  assign decB_fraction = _T_89[0:0]; // @[convert.scala 24:34]
  assign _T_92 = _T_63 == 1'h0; // @[convert.scala 25:26]
  assign _T_94 = _T_63 ? _T_81 : _T_80; // @[convert.scala 25:42]
  assign _T_97 = ~ _T_90; // @[convert.scala 26:67]
  assign _T_98 = _T_61 ? _T_97 : _T_90; // @[convert.scala 26:51]
  assign _T_99 = {_T_92,_T_94,_T_98}; // @[Cat.scala 29:58]
  assign _T_101 = io_B[3:0]; // @[convert.scala 29:56]
  assign _T_102 = _T_101 != 4'h0; // @[convert.scala 29:60]
  assign _T_103 = ~ _T_102; // @[convert.scala 29:41]
  assign decB_isNaR = _T_61 & _T_103; // @[convert.scala 29:39]
  assign _T_106 = _T_61 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_106 & _T_103; // @[convert.scala 30:41]
  assign _T_115 = realC[4]; // @[convert.scala 18:24]
  assign _T_116 = realC[3]; // @[convert.scala 18:40]
  assign _T_117 = _T_115 ^ _T_116; // @[convert.scala 18:36]
  assign _T_118 = realC[3:1]; // @[convert.scala 19:24]
  assign _T_119 = realC[2:0]; // @[convert.scala 19:43]
  assign _T_120 = _T_118 ^ _T_119; // @[convert.scala 19:39]
  assign _T_121 = _T_120[2:1]; // @[LZD.scala 43:32]
  assign _T_122 = _T_121 != 2'h0; // @[LZD.scala 39:14]
  assign _T_123 = _T_121[1]; // @[LZD.scala 39:21]
  assign _T_124 = _T_121[0]; // @[LZD.scala 39:30]
  assign _T_125 = ~ _T_124; // @[LZD.scala 39:27]
  assign _T_126 = _T_123 | _T_125; // @[LZD.scala 39:25]
  assign _T_127 = {_T_122,_T_126}; // @[Cat.scala 29:58]
  assign _T_128 = _T_120[0:0]; // @[LZD.scala 44:32]
  assign _T_130 = _T_127[1]; // @[Shift.scala 12:21]
  assign _T_132 = _T_127[0:0]; // @[LZD.scala 55:32]
  assign _T_133 = _T_130 ? _T_132 : _T_128; // @[LZD.scala 55:20]
  assign _T_134 = {_T_130,_T_133}; // @[Cat.scala 29:58]
  assign _T_135 = ~ _T_134; // @[convert.scala 21:22]
  assign _T_136 = realC[1:0]; // @[convert.scala 22:36]
  assign _T_137 = _T_135 < 2'h2; // @[Shift.scala 16:24]
  assign _T_138 = _T_135[0]; // @[Shift.scala 17:37]
  assign _T_140 = _T_136[0:0]; // @[Shift.scala 64:52]
  assign _T_141 = {_T_140,1'h0}; // @[Cat.scala 29:58]
  assign _T_142 = _T_138 ? _T_141 : _T_136; // @[Shift.scala 64:27]
  assign _T_143 = _T_137 ? _T_142 : 2'h0; // @[Shift.scala 16:10]
  assign _T_144 = _T_143[1:1]; // @[convert.scala 23:34]
  assign _T_146 = _T_117 == 1'h0; // @[convert.scala 25:26]
  assign _T_148 = _T_117 ? _T_135 : _T_134; // @[convert.scala 25:42]
  assign _T_151 = ~ _T_144; // @[convert.scala 26:67]
  assign _T_152 = _T_115 ? _T_151 : _T_144; // @[convert.scala 26:51]
  assign _T_153 = {_T_146,_T_148,_T_152}; // @[Cat.scala 29:58]
  assign _T_155 = realC[3:0]; // @[convert.scala 29:56]
  assign _T_156 = _T_155 != 4'h0; // @[convert.scala 29:60]
  assign _T_157 = ~ _T_156; // @[convert.scala 29:41]
  assign decC_isNaR = _T_115 & _T_157; // @[convert.scala 29:39]
  assign _T_160 = _T_115 == 1'h0; // @[convert.scala 30:19]
  assign _T_168 = decA_isNaR | decB_isNaR; // @[FMA_Dec.scala 46:30]
  assign _T_170 = ~ _T_7; // @[FMA_Dec.scala 49:34]
  assign _T_171 = ~ decA_isZero; // @[FMA_Dec.scala 49:47]
  assign _T_172 = _T_170 & _T_171; // @[FMA_Dec.scala 49:45]
  assign _T_174 = {_T_7,_T_172,decA_fraction}; // @[Cat.scala 29:58]
  assign _T_176 = ~ _T_61; // @[FMA_Dec.scala 50:34]
  assign _T_177 = ~ decB_isZero; // @[FMA_Dec.scala 50:47]
  assign _T_178 = _T_176 & _T_177; // @[FMA_Dec.scala 50:45]
  assign _T_180 = {_T_61,_T_178,decB_fraction}; // @[Cat.scala 29:58]
  assign io_sigA = $signed(_T_174); // @[FMA_Dec.scala 49:16]
  assign io_sigB = $signed(_T_180); // @[FMA_Dec.scala 50:16]
  assign io_outIsNaR = _T_168 | decC_isNaR; // @[FMA_Dec.scala 46:16]
  assign io_Csign = realC[4]; // @[FMA_Dec.scala 55:12]
  assign io_CisNar = _T_115 & _T_157; // @[FMA_Dec.scala 51:17]
  assign io_CisZero = _T_160 & _T_157; // @[FMA_Dec.scala 52:17]
  assign io_Cfrac = _T_143[0:0]; // @[FMA_Dec.scala 53:17]
  assign io_Ascale = $signed(_T_45); // @[FMA_Dec.scala 47:13]
  assign io_Bscale = $signed(_T_99); // @[FMA_Dec.scala 48:13]
  assign io_Cscale = $signed(_T_153); // @[FMA_Dec.scala 54:16]
endmodule
