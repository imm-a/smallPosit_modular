module PositDivSqrter7_1(
  input        clock,
  input        reset,
  output       io_inReady,
  input        io_inValid,
  input        io_sqrtOp,
  input  [6:0] io_A,
  input  [6:0] io_B,
  output       io_diviValid,
  output       io_sqrtValid,
  output       io_invalidExc,
  output [6:0] io_Q
);
  reg [3:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [5:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg [2:0] fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [9:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [9:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [4:0] _T_4; // @[convert.scala 19:24]
  wire [4:0] _T_5; // @[convert.scala 19:43]
  wire [4:0] _T_6; // @[convert.scala 19:39]
  wire [3:0] _T_7; // @[LZD.scala 43:32]
  wire [1:0] _T_8; // @[LZD.scala 43:32]
  wire  _T_9; // @[LZD.scala 39:14]
  wire  _T_10; // @[LZD.scala 39:21]
  wire  _T_11; // @[LZD.scala 39:30]
  wire  _T_12; // @[LZD.scala 39:27]
  wire  _T_13; // @[LZD.scala 39:25]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [1:0] _T_15; // @[LZD.scala 44:32]
  wire  _T_16; // @[LZD.scala 39:14]
  wire  _T_17; // @[LZD.scala 39:21]
  wire  _T_18; // @[LZD.scala 39:30]
  wire  _T_19; // @[LZD.scala 39:27]
  wire  _T_20; // @[LZD.scala 39:25]
  wire [1:0] _T_21; // @[Cat.scala 29:58]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[LZD.scala 49:16]
  wire  _T_25; // @[LZD.scala 49:27]
  wire  _T_26; // @[LZD.scala 49:25]
  wire  _T_27; // @[LZD.scala 49:47]
  wire  _T_28; // @[LZD.scala 49:59]
  wire  _T_29; // @[LZD.scala 49:35]
  wire [2:0] _T_31; // @[Cat.scala 29:58]
  wire  _T_32; // @[LZD.scala 44:32]
  wire  _T_34; // @[Shift.scala 12:21]
  wire [1:0] _T_36; // @[Cat.scala 29:58]
  wire [1:0] _T_37; // @[LZD.scala 55:32]
  wire [1:0] _T_38; // @[LZD.scala 55:20]
  wire [2:0] _T_39; // @[Cat.scala 29:58]
  wire [2:0] _T_40; // @[convert.scala 21:22]
  wire [3:0] _T_41; // @[convert.scala 22:36]
  wire  _T_42; // @[Shift.scala 16:24]
  wire [1:0] _T_43; // @[Shift.scala 17:37]
  wire  _T_44; // @[Shift.scala 12:21]
  wire [1:0] _T_45; // @[Shift.scala 64:52]
  wire [3:0] _T_47; // @[Cat.scala 29:58]
  wire [3:0] _T_48; // @[Shift.scala 64:27]
  wire  _T_49; // @[Shift.scala 66:70]
  wire [2:0] _T_51; // @[Shift.scala 64:52]
  wire [3:0] _T_52; // @[Cat.scala 29:58]
  wire [3:0] _T_53; // @[Shift.scala 64:27]
  wire [3:0] _T_54; // @[Shift.scala 16:10]
  wire  _T_55; // @[convert.scala 23:34]
  wire [2:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_57; // @[convert.scala 25:26]
  wire [2:0] _T_59; // @[convert.scala 25:42]
  wire  _T_62; // @[convert.scala 26:67]
  wire  _T_63; // @[convert.scala 26:51]
  wire [4:0] _T_64; // @[Cat.scala 29:58]
  wire [5:0] _T_66; // @[convert.scala 29:56]
  wire  _T_67; // @[convert.scala 29:60]
  wire  _T_68; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_71; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [4:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_80; // @[convert.scala 18:24]
  wire  _T_81; // @[convert.scala 18:40]
  wire  _T_82; // @[convert.scala 18:36]
  wire [4:0] _T_83; // @[convert.scala 19:24]
  wire [4:0] _T_84; // @[convert.scala 19:43]
  wire [4:0] _T_85; // @[convert.scala 19:39]
  wire [3:0] _T_86; // @[LZD.scala 43:32]
  wire [1:0] _T_87; // @[LZD.scala 43:32]
  wire  _T_88; // @[LZD.scala 39:14]
  wire  _T_89; // @[LZD.scala 39:21]
  wire  _T_90; // @[LZD.scala 39:30]
  wire  _T_91; // @[LZD.scala 39:27]
  wire  _T_92; // @[LZD.scala 39:25]
  wire [1:0] _T_93; // @[Cat.scala 29:58]
  wire [1:0] _T_94; // @[LZD.scala 44:32]
  wire  _T_95; // @[LZD.scala 39:14]
  wire  _T_96; // @[LZD.scala 39:21]
  wire  _T_97; // @[LZD.scala 39:30]
  wire  _T_98; // @[LZD.scala 39:27]
  wire  _T_99; // @[LZD.scala 39:25]
  wire [1:0] _T_100; // @[Cat.scala 29:58]
  wire  _T_101; // @[Shift.scala 12:21]
  wire  _T_102; // @[Shift.scala 12:21]
  wire  _T_103; // @[LZD.scala 49:16]
  wire  _T_104; // @[LZD.scala 49:27]
  wire  _T_105; // @[LZD.scala 49:25]
  wire  _T_106; // @[LZD.scala 49:47]
  wire  _T_107; // @[LZD.scala 49:59]
  wire  _T_108; // @[LZD.scala 49:35]
  wire [2:0] _T_110; // @[Cat.scala 29:58]
  wire  _T_111; // @[LZD.scala 44:32]
  wire  _T_113; // @[Shift.scala 12:21]
  wire [1:0] _T_115; // @[Cat.scala 29:58]
  wire [1:0] _T_116; // @[LZD.scala 55:32]
  wire [1:0] _T_117; // @[LZD.scala 55:20]
  wire [2:0] _T_118; // @[Cat.scala 29:58]
  wire [2:0] _T_119; // @[convert.scala 21:22]
  wire [3:0] _T_120; // @[convert.scala 22:36]
  wire  _T_121; // @[Shift.scala 16:24]
  wire [1:0] _T_122; // @[Shift.scala 17:37]
  wire  _T_123; // @[Shift.scala 12:21]
  wire [1:0] _T_124; // @[Shift.scala 64:52]
  wire [3:0] _T_126; // @[Cat.scala 29:58]
  wire [3:0] _T_127; // @[Shift.scala 64:27]
  wire  _T_128; // @[Shift.scala 66:70]
  wire [2:0] _T_130; // @[Shift.scala 64:52]
  wire [3:0] _T_131; // @[Cat.scala 29:58]
  wire [3:0] _T_132; // @[Shift.scala 64:27]
  wire [3:0] _T_133; // @[Shift.scala 16:10]
  wire  _T_134; // @[convert.scala 23:34]
  wire [2:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_136; // @[convert.scala 25:26]
  wire [2:0] _T_138; // @[convert.scala 25:42]
  wire  _T_141; // @[convert.scala 26:67]
  wire  _T_142; // @[convert.scala 26:51]
  wire [4:0] _T_143; // @[Cat.scala 29:58]
  wire [5:0] _T_145; // @[convert.scala 29:56]
  wire  _T_146; // @[convert.scala 29:60]
  wire  _T_147; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_150; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [4:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_159; // @[Bitwise.scala 71:12]
  wire  _T_160; // @[PositDivisionSqrt.scala 80:40]
  wire [9:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_163; // @[PositDivisionSqrt.scala 82:31]
  wire [9:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_166; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_167; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_168; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_169; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_170; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_171; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_172; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_173; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_174; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_175; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [5:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_178; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_179; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_180; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_181; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_182; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_183; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_184; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_185; // @[PositDivisionSqrt.scala 117:30]
  wire [3:0] _T_187; // @[PositDivisionSqrt.scala 119:26]
  wire [3:0] _T_188; // @[PositDivisionSqrt.scala 118:20]
  wire [3:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [3:0] _T_189; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_191; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_192; // @[PositDivisionSqrt.scala 123:27]
  wire [3:0] _T_194; // @[PositDivisionSqrt.scala 123:52]
  wire [3:0] _T_195; // @[PositDivisionSqrt.scala 123:20]
  wire [3:0] _T_196; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_198; // @[PositDivisionSqrt.scala 124:27]
  wire [3:0] _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _T_200; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _T_201; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_203; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_204; // @[PositDivisionSqrt.scala 137:28]
  wire [15:0] _T_205; // @[PositDivisionSqrt.scala 146:22]
  wire [13:0] _T_206; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_207; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_208; // @[PositDivisionSqrt.scala 148:23]
  wire [9:0] _T_209; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_210; // @[PositDivisionSqrt.scala 149:23]
  wire [10:0] _T_211; // @[PositDivisionSqrt.scala 149:46]
  wire [9:0] _T_212; // @[PositDivisionSqrt.scala 149:56]
  wire [9:0] _T_213; // @[PositDivisionSqrt.scala 149:16]
  wire [9:0] _T_214; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_215; // @[PositDivisionSqrt.scala 150:17]
  wire [9:0] _T_216; // @[PositDivisionSqrt.scala 150:16]
  wire [9:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_218; // @[PositDivisionSqrt.scala 152:29]
  wire [9:0] _T_219; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_220; // @[PositDivisionSqrt.scala 153:29]
  wire [6:0] _T_221; // @[PositDivisionSqrt.scala 153:22]
  wire [9:0] _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  wire [9:0] _T_222; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_224; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_225; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_226; // @[PositDivisionSqrt.scala 154:57]
  wire [9:0] _T_229; // @[Cat.scala 29:58]
  wire [9:0] _T_230; // @[PositDivisionSqrt.scala 154:22]
  wire [9:0] _T_231; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_233; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_234; // @[PositDivisionSqrt.scala 156:83]
  wire [5:0] _T_236; // @[Bitwise.scala 71:12]
  wire [8:0] bitMask; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  wire [8:0] _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  wire [8:0] _T_237; // @[PositDivisionSqrt.scala 156:53]
  wire [9:0] _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  wire [9:0] _T_238; // @[PositDivisionSqrt.scala 155:51]
  wire [7:0] _T_239; // @[PositDivisionSqrt.scala 157:53]
  wire [9:0] _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  wire [9:0] _T_240; // @[PositDivisionSqrt.scala 156:89]
  wire [9:0] _T_241; // @[PositDivisionSqrt.scala 155:22]
  wire [9:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_243; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_244; // @[PositDivisionSqrt.scala 162:40]
  wire [9:0] _T_247; // @[PositDivisionSqrt.scala 163:97]
  wire [9:0] _T_249; // @[PositDivisionSqrt.scala 164:97]
  wire [9:0] _T_250; // @[PositDivisionSqrt.scala 161:92]
  wire [10:0] _T_255; // @[PositDivisionSqrt.scala 168:98]
  wire [9:0] _T_256; // @[PositDivisionSqrt.scala 168:108]
  wire [9:0] _T_258; // @[PositDivisionSqrt.scala 168:112]
  wire [9:0] _T_262; // @[PositDivisionSqrt.scala 169:112]
  wire [9:0] _T_263; // @[PositDivisionSqrt.scala 166:26]
  wire [9:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_264; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_265; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_267; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_268; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_269; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_270; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_271; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_273; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_274; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_275; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_276; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_277; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_280; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_281; // @[PositDivisionSqrt.scala 187:28]
  wire [9:0] _T_284; // @[PositDivisionSqrt.scala 188:47]
  wire [9:0] _T_285; // @[PositDivisionSqrt.scala 188:18]
  wire [7:0] _T_287; // @[PositDivisionSqrt.scala 189:18]
  wire [9:0] _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  wire [9:0] _T_288; // @[PositDivisionSqrt.scala 188:78]
  wire [9:0] _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  wire [9:0] _T_290; // @[PositDivisionSqrt.scala 190:47]
  wire [9:0] _T_291; // @[PositDivisionSqrt.scala 190:18]
  wire [9:0] _T_292; // @[PositDivisionSqrt.scala 189:78]
  wire [1:0] _T_294; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [9:0] _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  wire [9:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire [2:0] _T_297; // @[PositDivisionSqrt.scala 200:97]
  wire [2:0] _T_298; // @[PositDivisionSqrt.scala 201:97]
  wire [2:0] realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_299; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_300; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_301; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  _T_303; // @[PositDivisionSqrt.scala 206:56]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_304; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_305; // @[Cat.scala 29:58]
  wire [2:0] _T_306; // @[PositDivisionSqrt.scala 209:63]
  wire [5:0] _GEN_18; // @[PositDivisionSqrt.scala 209:31]
  wire [5:0] _T_308; // @[PositDivisionSqrt.scala 209:31]
  wire [5:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [5:0] _T_310; // @[Mux.scala 87:16]
  wire [5:0] _T_311; // @[Mux.scala 87:16]
  wire [2:0] _T_312; // @[PositDivisionSqrt.scala 224:48]
  wire [2:0] _T_313; // @[PositDivisionSqrt.scala 224:64]
  wire [2:0] decQ_grs; // @[PositDivisionSqrt.scala 224:23]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [4:0] _GEN_19; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [4:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire  _T_319; // @[convert.scala 46:61]
  wire  _T_320; // @[convert.scala 46:52]
  wire  _T_322; // @[convert.scala 46:42]
  wire [3:0] _T_323; // @[convert.scala 48:34]
  wire  _T_324; // @[convert.scala 49:36]
  wire [3:0] _T_326; // @[convert.scala 50:36]
  wire [3:0] _T_327; // @[convert.scala 50:36]
  wire [3:0] _T_328; // @[convert.scala 50:28]
  wire  _T_329; // @[convert.scala 51:31]
  wire  _T_330; // @[convert.scala 52:43]
  wire [8:0] _T_334; // @[Cat.scala 29:58]
  wire [3:0] _T_335; // @[Shift.scala 39:17]
  wire  _T_336; // @[Shift.scala 39:24]
  wire  _T_338; // @[Shift.scala 90:30]
  wire [7:0] _T_339; // @[Shift.scala 90:48]
  wire  _T_340; // @[Shift.scala 90:57]
  wire  _T_341; // @[Shift.scala 90:39]
  wire  _T_342; // @[Shift.scala 12:21]
  wire  _T_343; // @[Shift.scala 12:21]
  wire [7:0] _T_345; // @[Bitwise.scala 71:12]
  wire [8:0] _T_346; // @[Cat.scala 29:58]
  wire [8:0] _T_347; // @[Shift.scala 91:22]
  wire [2:0] _T_348; // @[Shift.scala 92:77]
  wire [4:0] _T_349; // @[Shift.scala 90:30]
  wire [3:0] _T_350; // @[Shift.scala 90:48]
  wire  _T_351; // @[Shift.scala 90:57]
  wire [4:0] _GEN_20; // @[Shift.scala 90:39]
  wire [4:0] _T_352; // @[Shift.scala 90:39]
  wire  _T_353; // @[Shift.scala 12:21]
  wire  _T_354; // @[Shift.scala 12:21]
  wire [3:0] _T_356; // @[Bitwise.scala 71:12]
  wire [8:0] _T_357; // @[Cat.scala 29:58]
  wire [8:0] _T_358; // @[Shift.scala 91:22]
  wire [1:0] _T_359; // @[Shift.scala 92:77]
  wire [6:0] _T_360; // @[Shift.scala 90:30]
  wire [1:0] _T_361; // @[Shift.scala 90:48]
  wire  _T_362; // @[Shift.scala 90:57]
  wire [6:0] _GEN_21; // @[Shift.scala 90:39]
  wire [6:0] _T_363; // @[Shift.scala 90:39]
  wire  _T_364; // @[Shift.scala 12:21]
  wire  _T_365; // @[Shift.scala 12:21]
  wire [1:0] _T_367; // @[Bitwise.scala 71:12]
  wire [8:0] _T_368; // @[Cat.scala 29:58]
  wire [8:0] _T_369; // @[Shift.scala 91:22]
  wire  _T_370; // @[Shift.scala 92:77]
  wire [7:0] _T_371; // @[Shift.scala 90:30]
  wire  _T_372; // @[Shift.scala 90:48]
  wire [7:0] _GEN_22; // @[Shift.scala 90:39]
  wire [7:0] _T_374; // @[Shift.scala 90:39]
  wire  _T_376; // @[Shift.scala 12:21]
  wire [8:0] _T_377; // @[Cat.scala 29:58]
  wire [8:0] _T_378; // @[Shift.scala 91:22]
  wire [8:0] _T_381; // @[Bitwise.scala 71:12]
  wire [8:0] _T_382; // @[Shift.scala 39:10]
  wire  _T_383; // @[convert.scala 55:31]
  wire  _T_384; // @[convert.scala 56:31]
  wire  _T_385; // @[convert.scala 57:31]
  wire  _T_386; // @[convert.scala 58:31]
  wire [5:0] _T_387; // @[convert.scala 59:69]
  wire  _T_388; // @[convert.scala 59:81]
  wire  _T_389; // @[convert.scala 59:50]
  wire  _T_391; // @[convert.scala 60:81]
  wire  _T_392; // @[convert.scala 61:44]
  wire  _T_393; // @[convert.scala 61:52]
  wire  _T_394; // @[convert.scala 61:36]
  wire  _T_395; // @[convert.scala 62:63]
  wire  _T_396; // @[convert.scala 62:103]
  wire  _T_397; // @[convert.scala 62:60]
  wire [5:0] _GEN_23; // @[convert.scala 63:56]
  wire [5:0] _T_400; // @[convert.scala 63:56]
  wire [6:0] _T_401; // @[Cat.scala 29:58]
  wire [6:0] _T_403; // @[Mux.scala 87:16]
  assign _T_1 = io_A[6]; // @[convert.scala 18:24]
  assign _T_2 = io_A[5]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[5:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[4:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[4:1]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[3:2]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8 != 2'h0; // @[LZD.scala 39:14]
  assign _T_10 = _T_8[1]; // @[LZD.scala 39:21]
  assign _T_11 = _T_8[0]; // @[LZD.scala 39:30]
  assign _T_12 = ~ _T_11; // @[LZD.scala 39:27]
  assign _T_13 = _T_10 | _T_12; // @[LZD.scala 39:25]
  assign _T_14 = {_T_9,_T_13}; // @[Cat.scala 29:58]
  assign _T_15 = _T_7[1:0]; // @[LZD.scala 44:32]
  assign _T_16 = _T_15 != 2'h0; // @[LZD.scala 39:14]
  assign _T_17 = _T_15[1]; // @[LZD.scala 39:21]
  assign _T_18 = _T_15[0]; // @[LZD.scala 39:30]
  assign _T_19 = ~ _T_18; // @[LZD.scala 39:27]
  assign _T_20 = _T_17 | _T_19; // @[LZD.scala 39:25]
  assign _T_21 = {_T_16,_T_20}; // @[Cat.scala 29:58]
  assign _T_22 = _T_14[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22 | _T_23; // @[LZD.scala 49:16]
  assign _T_25 = ~ _T_23; // @[LZD.scala 49:27]
  assign _T_26 = _T_22 | _T_25; // @[LZD.scala 49:25]
  assign _T_27 = _T_14[0:0]; // @[LZD.scala 49:47]
  assign _T_28 = _T_21[0:0]; // @[LZD.scala 49:59]
  assign _T_29 = _T_22 ? _T_27 : _T_28; // @[LZD.scala 49:35]
  assign _T_31 = {_T_24,_T_26,_T_29}; // @[Cat.scala 29:58]
  assign _T_32 = _T_6[0:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_31[2]; // @[Shift.scala 12:21]
  assign _T_36 = {1'h1,_T_32}; // @[Cat.scala 29:58]
  assign _T_37 = _T_31[1:0]; // @[LZD.scala 55:32]
  assign _T_38 = _T_34 ? _T_37 : _T_36; // @[LZD.scala 55:20]
  assign _T_39 = {_T_34,_T_38}; // @[Cat.scala 29:58]
  assign _T_40 = ~ _T_39; // @[convert.scala 21:22]
  assign _T_41 = io_A[3:0]; // @[convert.scala 22:36]
  assign _T_42 = _T_40 < 3'h4; // @[Shift.scala 16:24]
  assign _T_43 = _T_40[1:0]; // @[Shift.scala 17:37]
  assign _T_44 = _T_43[1]; // @[Shift.scala 12:21]
  assign _T_45 = _T_41[1:0]; // @[Shift.scala 64:52]
  assign _T_47 = {_T_45,2'h0}; // @[Cat.scala 29:58]
  assign _T_48 = _T_44 ? _T_47 : _T_41; // @[Shift.scala 64:27]
  assign _T_49 = _T_43[0:0]; // @[Shift.scala 66:70]
  assign _T_51 = _T_48[2:0]; // @[Shift.scala 64:52]
  assign _T_52 = {_T_51,1'h0}; // @[Cat.scala 29:58]
  assign _T_53 = _T_49 ? _T_52 : _T_48; // @[Shift.scala 64:27]
  assign _T_54 = _T_42 ? _T_53 : 4'h0; // @[Shift.scala 16:10]
  assign _T_55 = _T_54[3:3]; // @[convert.scala 23:34]
  assign decA_fraction = _T_54[2:0]; // @[convert.scala 24:34]
  assign _T_57 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_59 = _T_3 ? _T_40 : _T_39; // @[convert.scala 25:42]
  assign _T_62 = ~ _T_55; // @[convert.scala 26:67]
  assign _T_63 = _T_1 ? _T_62 : _T_55; // @[convert.scala 26:51]
  assign _T_64 = {_T_57,_T_59,_T_63}; // @[Cat.scala 29:58]
  assign _T_66 = io_A[5:0]; // @[convert.scala 29:56]
  assign _T_67 = _T_66 != 6'h0; // @[convert.scala 29:60]
  assign _T_68 = ~ _T_67; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_68; // @[convert.scala 29:39]
  assign _T_71 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_71 & _T_68; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_64); // @[convert.scala 32:24]
  assign _T_80 = io_B[6]; // @[convert.scala 18:24]
  assign _T_81 = io_B[5]; // @[convert.scala 18:40]
  assign _T_82 = _T_80 ^ _T_81; // @[convert.scala 18:36]
  assign _T_83 = io_B[5:1]; // @[convert.scala 19:24]
  assign _T_84 = io_B[4:0]; // @[convert.scala 19:43]
  assign _T_85 = _T_83 ^ _T_84; // @[convert.scala 19:39]
  assign _T_86 = _T_85[4:1]; // @[LZD.scala 43:32]
  assign _T_87 = _T_86[3:2]; // @[LZD.scala 43:32]
  assign _T_88 = _T_87 != 2'h0; // @[LZD.scala 39:14]
  assign _T_89 = _T_87[1]; // @[LZD.scala 39:21]
  assign _T_90 = _T_87[0]; // @[LZD.scala 39:30]
  assign _T_91 = ~ _T_90; // @[LZD.scala 39:27]
  assign _T_92 = _T_89 | _T_91; // @[LZD.scala 39:25]
  assign _T_93 = {_T_88,_T_92}; // @[Cat.scala 29:58]
  assign _T_94 = _T_86[1:0]; // @[LZD.scala 44:32]
  assign _T_95 = _T_94 != 2'h0; // @[LZD.scala 39:14]
  assign _T_96 = _T_94[1]; // @[LZD.scala 39:21]
  assign _T_97 = _T_94[0]; // @[LZD.scala 39:30]
  assign _T_98 = ~ _T_97; // @[LZD.scala 39:27]
  assign _T_99 = _T_96 | _T_98; // @[LZD.scala 39:25]
  assign _T_100 = {_T_95,_T_99}; // @[Cat.scala 29:58]
  assign _T_101 = _T_93[1]; // @[Shift.scala 12:21]
  assign _T_102 = _T_100[1]; // @[Shift.scala 12:21]
  assign _T_103 = _T_101 | _T_102; // @[LZD.scala 49:16]
  assign _T_104 = ~ _T_102; // @[LZD.scala 49:27]
  assign _T_105 = _T_101 | _T_104; // @[LZD.scala 49:25]
  assign _T_106 = _T_93[0:0]; // @[LZD.scala 49:47]
  assign _T_107 = _T_100[0:0]; // @[LZD.scala 49:59]
  assign _T_108 = _T_101 ? _T_106 : _T_107; // @[LZD.scala 49:35]
  assign _T_110 = {_T_103,_T_105,_T_108}; // @[Cat.scala 29:58]
  assign _T_111 = _T_85[0:0]; // @[LZD.scala 44:32]
  assign _T_113 = _T_110[2]; // @[Shift.scala 12:21]
  assign _T_115 = {1'h1,_T_111}; // @[Cat.scala 29:58]
  assign _T_116 = _T_110[1:0]; // @[LZD.scala 55:32]
  assign _T_117 = _T_113 ? _T_116 : _T_115; // @[LZD.scala 55:20]
  assign _T_118 = {_T_113,_T_117}; // @[Cat.scala 29:58]
  assign _T_119 = ~ _T_118; // @[convert.scala 21:22]
  assign _T_120 = io_B[3:0]; // @[convert.scala 22:36]
  assign _T_121 = _T_119 < 3'h4; // @[Shift.scala 16:24]
  assign _T_122 = _T_119[1:0]; // @[Shift.scala 17:37]
  assign _T_123 = _T_122[1]; // @[Shift.scala 12:21]
  assign _T_124 = _T_120[1:0]; // @[Shift.scala 64:52]
  assign _T_126 = {_T_124,2'h0}; // @[Cat.scala 29:58]
  assign _T_127 = _T_123 ? _T_126 : _T_120; // @[Shift.scala 64:27]
  assign _T_128 = _T_122[0:0]; // @[Shift.scala 66:70]
  assign _T_130 = _T_127[2:0]; // @[Shift.scala 64:52]
  assign _T_131 = {_T_130,1'h0}; // @[Cat.scala 29:58]
  assign _T_132 = _T_128 ? _T_131 : _T_127; // @[Shift.scala 64:27]
  assign _T_133 = _T_121 ? _T_132 : 4'h0; // @[Shift.scala 16:10]
  assign _T_134 = _T_133[3:3]; // @[convert.scala 23:34]
  assign decB_fraction = _T_133[2:0]; // @[convert.scala 24:34]
  assign _T_136 = _T_82 == 1'h0; // @[convert.scala 25:26]
  assign _T_138 = _T_82 ? _T_119 : _T_118; // @[convert.scala 25:42]
  assign _T_141 = ~ _T_134; // @[convert.scala 26:67]
  assign _T_142 = _T_80 ? _T_141 : _T_134; // @[convert.scala 26:51]
  assign _T_143 = {_T_136,_T_138,_T_142}; // @[Cat.scala 29:58]
  assign _T_145 = io_B[5:0]; // @[convert.scala 29:56]
  assign _T_146 = _T_145 != 6'h0; // @[convert.scala 29:60]
  assign _T_147 = ~ _T_146; // @[convert.scala 29:41]
  assign decB_isNaR = _T_80 & _T_147; // @[convert.scala 29:39]
  assign _T_150 = _T_80 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_150 & _T_147; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_143); // @[convert.scala 32:24]
  assign _T_159 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_160 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_159,_T_160,decA_fraction,3'h0}; // @[Cat.scala 29:58]
  assign _T_163 = ~ _T_80; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_80,_T_163,decB_fraction,5'h0}; // @[Cat.scala 29:58]
  assign _T_166 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_166 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_167 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_168 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_169 = _T_168 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_170 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_171 = decA_isZero & _T_170; // @[PositDivisionSqrt.scala 94:43]
  assign _T_172 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_173 = _T_171 & _T_172; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_174 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_175 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_174 & _T_175; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_174 & _T_71; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_178 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_178; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 4'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_179 = sigX_Z[9]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_180 = sigX_Z[7]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_179 ^ _T_180; // @[PositDivisionSqrt.scala 113:50]
  assign _T_181 = cycleNum == 4'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_181 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_182 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_183 = _T_182 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_184 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_185 = entering & _T_184; // @[PositDivisionSqrt.scala 117:30]
  assign _T_187 = io_sqrtOp ? 4'h8 : 4'ha; // @[PositDivisionSqrt.scala 119:26]
  assign _T_188 = entering_normalCase ? _T_187 : 4'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{3'd0}, _T_185}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_189 = _GEN_9 | _T_188; // @[PositDivisionSqrt.scala 117:64]
  assign _T_191 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_192 = _T_182 & _T_191; // @[PositDivisionSqrt.scala 123:27]
  assign _T_194 = cycleNum - 4'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_195 = _T_192 ? _T_194 : 4'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _T_196 = _T_189 | _T_195; // @[PositDivisionSqrt.scala 122:64]
  assign _T_198 = _T_182 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_10 = {{3'd0}, _T_198}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_200 = _T_196 | _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  assign _T_201 = decA_scale[4:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_203 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_204 = entering_normalCase & _T_203; // @[PositDivisionSqrt.scala 137:28]
  assign _T_205 = 16'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign _T_206 = _T_205[15:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_207 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_208 = ready & _T_207; // @[PositDivisionSqrt.scala 148:23]
  assign _T_209 = _T_208 ? sigA_S : 10'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_210 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_211 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_212 = _T_211[9:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_213 = _T_210 ? _T_212 : 10'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_214 = _T_209 | _T_213; // @[PositDivisionSqrt.scala 148:66]
  assign _T_215 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_216 = _T_215 ? rem_Z : 10'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_214 | _T_216; // @[PositDivisionSqrt.scala 149:66]
  assign _T_218 = ready & _T_203; // @[PositDivisionSqrt.scala 152:29]
  assign _T_219 = _T_218 ? sigB_S : 10'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_220 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_221 = _T_220 ? 7'h40 : 7'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_11 = {{3'd0}, _T_221}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_222 = _T_219 | _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  assign _T_224 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_225 = _T_215 & _T_224; // @[PositDivisionSqrt.scala 154:30]
  assign _T_226 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_229 = {signB_Z,_T_226,fractB_Z,5'h0}; // @[Cat.scala 29:58]
  assign _T_230 = _T_225 ? _T_229 : 10'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_231 = _T_222 | _T_230; // @[PositDivisionSqrt.scala 153:93]
  assign _T_233 = _T_215 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_234 = rem[9:9]; // @[PositDivisionSqrt.scala 156:83]
  assign _T_236 = _T_234 ? 6'h3f : 6'h0; // @[Bitwise.scala 71:12]
  assign bitMask = _T_206[8:0]; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  assign _GEN_12 = {{3'd0}, _T_236}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_237 = bitMask & _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_13 = {{1'd0}, _T_237}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_238 = sigX_Z | _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  assign _T_239 = bitMask[8:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_14 = {{2'd0}, _T_239}; // @[PositDivisionSqrt.scala 156:89]
  assign _T_240 = _T_238 | _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  assign _T_241 = _T_233 ? _T_240 : 10'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_231 | _T_241; // @[PositDivisionSqrt.scala 154:93]
  assign _T_243 = trialTerm[9:9]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_244 = _T_234 ^ _T_243; // @[PositDivisionSqrt.scala 162:40]
  assign _T_247 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_249 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_250 = _T_244 ? _T_247 : _T_249; // @[PositDivisionSqrt.scala 161:92]
  assign _T_255 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_256 = _T_255[9:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_258 = _T_256 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_262 = _T_256 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_263 = _T_244 ? _T_258 : _T_262; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_250 : _T_263; // @[PositDivisionSqrt.scala 159:27]
  assign _T_264 = trialRem != 10'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_264 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_265 = rem != 10'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_265 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_267 = trialRem[9:9]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_268 = _T_243 ^ _T_267; // @[PositDivisionSqrt.scala 176:49]
  assign _T_269 = ~ _T_268; // @[PositDivisionSqrt.scala 176:29]
  assign _T_270 = sigX_Z[9:9]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_271 = ~ _T_270; // @[PositDivisionSqrt.scala 178:49]
  assign _T_273 = remIsZero ? _T_270 : _T_269; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_271 : _T_273; // @[Mux.scala 87:16]
  assign _T_274 = cycleNum > 4'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_275 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_276 = _T_274 & _T_275; // @[PositDivisionSqrt.scala 183:48]
  assign _T_277 = entering_normalCase | _T_276; // @[PositDivisionSqrt.scala 183:28]
  assign _T_280 = _T_215 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_281 = entering_normalCase | _T_280; // @[PositDivisionSqrt.scala 187:28]
  assign _T_284 = {newBit, 9'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_285 = _T_218 ? _T_284 : 10'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_287 = _T_220 ? 8'h80 : 8'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_15 = {{2'd0}, _T_287}; // @[PositDivisionSqrt.scala 188:78]
  assign _T_288 = _T_285 | _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  assign _GEN_16 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_290 = sigX_Z | _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  assign _T_291 = _T_215 ? _T_290 : 10'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_292 = _T_288 | _T_291; // @[PositDivisionSqrt.scala 189:78]
  assign _T_294 = {_T_270, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_294 : {{1'd0}, _T_270}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_17 = {{8'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  assign _T_297 = realSigX[6:4]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_298 = realSigX[5:3]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_297 : _T_298; // @[PositDivisionSqrt.scala 198:21]
  assign _T_299 = realSigX[9]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_300 = realSigX[7]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_301 = _T_299 ^ _T_300; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_301; // @[PositDivisionSqrt.scala 205:23]
  assign _T_303 = realSigX[6]; // @[PositDivisionSqrt.scala 206:56]
  assign notNeedSubTwo = _T_299 ^ _T_303; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_304 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_304; // @[PositDivisionSqrt.scala 208:36]
  assign _T_305 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_306 = {1'b0,$signed(_T_305)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_18 = {{3{_T_306[2]}},_T_306}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_308 = $signed(scale_Z) - $signed(_GEN_18); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_308); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-6'shb); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(6'sha); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[9:9]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_310 = underflow ? $signed(-6'shb) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_311 = overflow ? $signed(6'sha) : $signed(_T_310); // @[Mux.scala 87:16]
  assign _T_312 = realSigX[3:1]; // @[PositDivisionSqrt.scala 224:48]
  assign _T_313 = realSigX[2:0]; // @[PositDivisionSqrt.scala 224:64]
  assign decQ_grs = scaleNotChange ? _T_312 : _T_313; // @[PositDivisionSqrt.scala 224:23]
  assign outValid = cycleNum == 4'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_19 = _T_311[4:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_19); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_319 = decQ_scale[0]; // @[convert.scala 46:61]
  assign _T_320 = ~ _T_319; // @[convert.scala 46:52]
  assign _T_322 = decQ_sign ? _T_320 : _T_319; // @[convert.scala 46:42]
  assign _T_323 = decQ_scale[4:1]; // @[convert.scala 48:34]
  assign _T_324 = _T_323[3:3]; // @[convert.scala 49:36]
  assign _T_326 = ~ _T_323; // @[convert.scala 50:36]
  assign _T_327 = $signed(_T_326); // @[convert.scala 50:36]
  assign _T_328 = _T_324 ? $signed(_T_327) : $signed(_T_323); // @[convert.scala 50:28]
  assign _T_329 = _T_324 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_330 = ~ _T_329; // @[convert.scala 52:43]
  assign _T_334 = {_T_330,_T_329,_T_322,realFrac,decQ_grs}; // @[Cat.scala 29:58]
  assign _T_335 = $unsigned(_T_328); // @[Shift.scala 39:17]
  assign _T_336 = _T_335 < 4'h9; // @[Shift.scala 39:24]
  assign _T_338 = _T_334[8:8]; // @[Shift.scala 90:30]
  assign _T_339 = _T_334[7:0]; // @[Shift.scala 90:48]
  assign _T_340 = _T_339 != 8'h0; // @[Shift.scala 90:57]
  assign _T_341 = _T_338 | _T_340; // @[Shift.scala 90:39]
  assign _T_342 = _T_335[3]; // @[Shift.scala 12:21]
  assign _T_343 = _T_334[8]; // @[Shift.scala 12:21]
  assign _T_345 = _T_343 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_346 = {_T_345,_T_341}; // @[Cat.scala 29:58]
  assign _T_347 = _T_342 ? _T_346 : _T_334; // @[Shift.scala 91:22]
  assign _T_348 = _T_335[2:0]; // @[Shift.scala 92:77]
  assign _T_349 = _T_347[8:4]; // @[Shift.scala 90:30]
  assign _T_350 = _T_347[3:0]; // @[Shift.scala 90:48]
  assign _T_351 = _T_350 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{4'd0}, _T_351}; // @[Shift.scala 90:39]
  assign _T_352 = _T_349 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_353 = _T_348[2]; // @[Shift.scala 12:21]
  assign _T_354 = _T_347[8]; // @[Shift.scala 12:21]
  assign _T_356 = _T_354 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_357 = {_T_356,_T_352}; // @[Cat.scala 29:58]
  assign _T_358 = _T_353 ? _T_357 : _T_347; // @[Shift.scala 91:22]
  assign _T_359 = _T_348[1:0]; // @[Shift.scala 92:77]
  assign _T_360 = _T_358[8:2]; // @[Shift.scala 90:30]
  assign _T_361 = _T_358[1:0]; // @[Shift.scala 90:48]
  assign _T_362 = _T_361 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{6'd0}, _T_362}; // @[Shift.scala 90:39]
  assign _T_363 = _T_360 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_364 = _T_359[1]; // @[Shift.scala 12:21]
  assign _T_365 = _T_358[8]; // @[Shift.scala 12:21]
  assign _T_367 = _T_365 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_368 = {_T_367,_T_363}; // @[Cat.scala 29:58]
  assign _T_369 = _T_364 ? _T_368 : _T_358; // @[Shift.scala 91:22]
  assign _T_370 = _T_359[0:0]; // @[Shift.scala 92:77]
  assign _T_371 = _T_369[8:1]; // @[Shift.scala 90:30]
  assign _T_372 = _T_369[0:0]; // @[Shift.scala 90:48]
  assign _GEN_22 = {{7'd0}, _T_372}; // @[Shift.scala 90:39]
  assign _T_374 = _T_371 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_376 = _T_369[8]; // @[Shift.scala 12:21]
  assign _T_377 = {_T_376,_T_374}; // @[Cat.scala 29:58]
  assign _T_378 = _T_370 ? _T_377 : _T_369; // @[Shift.scala 91:22]
  assign _T_381 = _T_343 ? 9'h1ff : 9'h0; // @[Bitwise.scala 71:12]
  assign _T_382 = _T_336 ? _T_378 : _T_381; // @[Shift.scala 39:10]
  assign _T_383 = _T_382[3]; // @[convert.scala 55:31]
  assign _T_384 = _T_382[2]; // @[convert.scala 56:31]
  assign _T_385 = _T_382[1]; // @[convert.scala 57:31]
  assign _T_386 = _T_382[0]; // @[convert.scala 58:31]
  assign _T_387 = _T_382[8:3]; // @[convert.scala 59:69]
  assign _T_388 = _T_387 != 6'h0; // @[convert.scala 59:81]
  assign _T_389 = ~ _T_388; // @[convert.scala 59:50]
  assign _T_391 = _T_387 == 6'h3f; // @[convert.scala 60:81]
  assign _T_392 = _T_383 | _T_385; // @[convert.scala 61:44]
  assign _T_393 = _T_392 | _T_386; // @[convert.scala 61:52]
  assign _T_394 = _T_384 & _T_393; // @[convert.scala 61:36]
  assign _T_395 = ~ _T_391; // @[convert.scala 62:63]
  assign _T_396 = _T_395 & _T_394; // @[convert.scala 62:103]
  assign _T_397 = _T_389 | _T_396; // @[convert.scala 62:60]
  assign _GEN_23 = {{5'd0}, _T_397}; // @[convert.scala 63:56]
  assign _T_400 = _T_387 + _GEN_23; // @[convert.scala 63:56]
  assign _T_401 = {decQ_sign,_T_400}; // @[Cat.scala 29:58]
  assign _T_403 = isZero_Z ? 7'h0 : _T_401; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_224; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 7'h40 : _T_403; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 4'h0;
    end else begin
      if (_T_183) begin
        cycleNum <= _T_200;
      end
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_167;
      end else begin
        isNaR_Z <= _T_169;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_173;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_201[3]}},_T_201};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_204) begin
      signB_Z <= _T_80;
    end
    if (_T_204) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_277) begin
      if (ready) begin
        if (_T_244) begin
          rem_Z <= _T_247;
        end else begin
          rem_Z <= _T_249;
        end
      end else begin
        if (_T_244) begin
          rem_Z <= _T_258;
        end else begin
          rem_Z <= _T_262;
        end
      end
    end
    if (_T_281) begin
      sigX_Z <= _T_292;
    end
  end
endmodule
