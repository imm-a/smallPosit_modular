module PositFMA5_0(
  input        clock,
  input        reset,
  input        io_inValid,
  input  [1:0] io_fmaOp,
  input  [4:0] io_A,
  input  [4:0] io_B,
  input  [4:0] io_C,
  output [4:0] io_F,
  output       io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [4:0] _T_2; // @[Bitwise.scala 71:12]
  wire [4:0] _T_3; // @[PositFMA.scala 47:41]
  wire [4:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [4:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [4:0] _T_8; // @[Bitwise.scala 71:12]
  wire [4:0] _T_9; // @[PositFMA.scala 48:41]
  wire [4:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [4:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [2:0] _T_16; // @[convert.scala 19:24]
  wire [2:0] _T_17; // @[convert.scala 19:43]
  wire [2:0] _T_18; // @[convert.scala 19:39]
  wire [1:0] _T_19; // @[LZD.scala 43:32]
  wire  _T_20; // @[LZD.scala 39:14]
  wire  _T_21; // @[LZD.scala 39:21]
  wire  _T_22; // @[LZD.scala 39:30]
  wire  _T_23; // @[LZD.scala 39:27]
  wire  _T_24; // @[LZD.scala 39:25]
  wire [1:0] _T_25; // @[Cat.scala 29:58]
  wire  _T_26; // @[LZD.scala 44:32]
  wire  _T_28; // @[Shift.scala 12:21]
  wire  _T_30; // @[LZD.scala 55:32]
  wire  _T_31; // @[LZD.scala 55:20]
  wire [1:0] _T_32; // @[Cat.scala 29:58]
  wire [1:0] _T_33; // @[convert.scala 21:22]
  wire [1:0] _T_34; // @[convert.scala 22:36]
  wire  _T_35; // @[Shift.scala 16:24]
  wire  _T_36; // @[Shift.scala 17:37]
  wire  _T_38; // @[Shift.scala 64:52]
  wire [1:0] _T_39; // @[Cat.scala 29:58]
  wire [1:0] _T_40; // @[Shift.scala 64:27]
  wire [1:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_44; // @[convert.scala 25:26]
  wire [1:0] _T_46; // @[convert.scala 25:42]
  wire [2:0] _T_47; // @[Cat.scala 29:58]
  wire [3:0] _T_49; // @[convert.scala 29:56]
  wire  _T_50; // @[convert.scala 29:60]
  wire  _T_51; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_54; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [2:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_63; // @[convert.scala 18:24]
  wire  _T_64; // @[convert.scala 18:40]
  wire  _T_65; // @[convert.scala 18:36]
  wire [2:0] _T_66; // @[convert.scala 19:24]
  wire [2:0] _T_67; // @[convert.scala 19:43]
  wire [2:0] _T_68; // @[convert.scala 19:39]
  wire [1:0] _T_69; // @[LZD.scala 43:32]
  wire  _T_70; // @[LZD.scala 39:14]
  wire  _T_71; // @[LZD.scala 39:21]
  wire  _T_72; // @[LZD.scala 39:30]
  wire  _T_73; // @[LZD.scala 39:27]
  wire  _T_74; // @[LZD.scala 39:25]
  wire [1:0] _T_75; // @[Cat.scala 29:58]
  wire  _T_76; // @[LZD.scala 44:32]
  wire  _T_78; // @[Shift.scala 12:21]
  wire  _T_80; // @[LZD.scala 55:32]
  wire  _T_81; // @[LZD.scala 55:20]
  wire [1:0] _T_82; // @[Cat.scala 29:58]
  wire [1:0] _T_83; // @[convert.scala 21:22]
  wire [1:0] _T_84; // @[convert.scala 22:36]
  wire  _T_85; // @[Shift.scala 16:24]
  wire  _T_86; // @[Shift.scala 17:37]
  wire  _T_88; // @[Shift.scala 64:52]
  wire [1:0] _T_89; // @[Cat.scala 29:58]
  wire [1:0] _T_90; // @[Shift.scala 64:27]
  wire [1:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_94; // @[convert.scala 25:26]
  wire [1:0] _T_96; // @[convert.scala 25:42]
  wire [2:0] _T_97; // @[Cat.scala 29:58]
  wire [3:0] _T_99; // @[convert.scala 29:56]
  wire  _T_100; // @[convert.scala 29:60]
  wire  _T_101; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_104; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [2:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_113; // @[convert.scala 18:24]
  wire  _T_114; // @[convert.scala 18:40]
  wire  _T_115; // @[convert.scala 18:36]
  wire [2:0] _T_116; // @[convert.scala 19:24]
  wire [2:0] _T_117; // @[convert.scala 19:43]
  wire [2:0] _T_118; // @[convert.scala 19:39]
  wire [1:0] _T_119; // @[LZD.scala 43:32]
  wire  _T_120; // @[LZD.scala 39:14]
  wire  _T_121; // @[LZD.scala 39:21]
  wire  _T_122; // @[LZD.scala 39:30]
  wire  _T_123; // @[LZD.scala 39:27]
  wire  _T_124; // @[LZD.scala 39:25]
  wire [1:0] _T_125; // @[Cat.scala 29:58]
  wire  _T_126; // @[LZD.scala 44:32]
  wire  _T_128; // @[Shift.scala 12:21]
  wire  _T_130; // @[LZD.scala 55:32]
  wire  _T_131; // @[LZD.scala 55:20]
  wire [1:0] _T_132; // @[Cat.scala 29:58]
  wire [1:0] _T_133; // @[convert.scala 21:22]
  wire [1:0] _T_134; // @[convert.scala 22:36]
  wire  _T_135; // @[Shift.scala 16:24]
  wire  _T_136; // @[Shift.scala 17:37]
  wire  _T_138; // @[Shift.scala 64:52]
  wire [1:0] _T_139; // @[Cat.scala 29:58]
  wire  _T_144; // @[convert.scala 25:26]
  wire [1:0] _T_146; // @[convert.scala 25:42]
  wire [2:0] _T_147; // @[Cat.scala 29:58]
  wire [3:0] _T_149; // @[convert.scala 29:56]
  wire  _T_150; // @[convert.scala 29:60]
  wire  _T_151; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_154; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [2:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_162; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_163; // @[PositFMA.scala 59:34]
  wire  _T_164; // @[PositFMA.scala 59:47]
  wire  _T_165; // @[PositFMA.scala 59:45]
  wire [3:0] _T_167; // @[Cat.scala 29:58]
  wire [3:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_168; // @[PositFMA.scala 60:34]
  wire  _T_169; // @[PositFMA.scala 60:47]
  wire  _T_170; // @[PositFMA.scala 60:45]
  wire [3:0] _T_172; // @[Cat.scala 29:58]
  wire [3:0] sigB; // @[PositFMA.scala 60:76]
  wire [7:0] _T_173; // @[PositFMA.scala 62:25]
  wire [7:0] sigP; // @[PositFMA.scala 62:33]
  wire [1:0] head2; // @[PositFMA.scala 63:28]
  wire  _T_174; // @[PositFMA.scala 64:31]
  wire  _T_175; // @[PositFMA.scala 64:25]
  wire  _T_176; // @[PositFMA.scala 64:42]
  wire  addTwo; // @[PositFMA.scala 64:35]
  wire  _T_177; // @[PositFMA.scala 66:23]
  wire  _T_178; // @[PositFMA.scala 66:49]
  wire  addOne; // @[PositFMA.scala 66:43]
  wire [1:0] _T_179; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 67:39]
  wire  mulSign; // @[PositFMA.scala 68:28]
  wire [3:0] _T_180; // @[PositFMA.scala 70:30]
  wire [3:0] _GEN_12; // @[PositFMA.scala 70:44]
  wire [3:0] _T_182; // @[PositFMA.scala 70:44]
  wire [3:0] mulScale; // @[PositFMA.scala 70:44]
  wire [5:0] _T_183; // @[PositFMA.scala 73:29]
  wire [4:0] _T_184; // @[PositFMA.scala 74:29]
  wire [5:0] _T_185; // @[PositFMA.scala 74:48]
  wire [5:0] mulSigTmp; // @[PositFMA.scala 71:22]
  wire  _T_187; // @[PositFMA.scala 78:39]
  wire  _T_188; // @[PositFMA.scala 78:43]
  wire [4:0] _T_189; // @[PositFMA.scala 79:39]
  wire [6:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [6:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [1:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [3:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [2:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_215; // @[PositFMA.scala 108:29]
  wire  _T_216; // @[PositFMA.scala 108:47]
  wire  _T_217; // @[PositFMA.scala 108:45]
  wire [6:0] extAddSig; // @[Cat.scala 29:58]
  wire [3:0] _GEN_13; // @[PositFMA.scala 112:39]
  wire  mulGreater; // @[PositFMA.scala 112:39]
  wire [3:0] greaterScale; // @[PositFMA.scala 113:26]
  wire [3:0] smallerScale; // @[PositFMA.scala 114:26]
  wire [3:0] _T_221; // @[PositFMA.scala 115:36]
  wire [3:0] scaleDiff; // @[PositFMA.scala 115:36]
  wire [6:0] greaterSig; // @[PositFMA.scala 116:26]
  wire [6:0] smallerSigTmp; // @[PositFMA.scala 117:26]
  wire [3:0] _T_222; // @[PositFMA.scala 118:69]
  wire  _T_223; // @[Shift.scala 39:24]
  wire [2:0] _T_224; // @[Shift.scala 40:44]
  wire [2:0] _T_225; // @[Shift.scala 90:30]
  wire [3:0] _T_226; // @[Shift.scala 90:48]
  wire  _T_227; // @[Shift.scala 90:57]
  wire [2:0] _GEN_14; // @[Shift.scala 90:39]
  wire [2:0] _T_228; // @[Shift.scala 90:39]
  wire  _T_229; // @[Shift.scala 12:21]
  wire  _T_230; // @[Shift.scala 12:21]
  wire [3:0] _T_232; // @[Bitwise.scala 71:12]
  wire [6:0] _T_233; // @[Cat.scala 29:58]
  wire [6:0] _T_234; // @[Shift.scala 91:22]
  wire [1:0] _T_235; // @[Shift.scala 92:77]
  wire [4:0] _T_236; // @[Shift.scala 90:30]
  wire [1:0] _T_237; // @[Shift.scala 90:48]
  wire  _T_238; // @[Shift.scala 90:57]
  wire [4:0] _GEN_15; // @[Shift.scala 90:39]
  wire [4:0] _T_239; // @[Shift.scala 90:39]
  wire  _T_240; // @[Shift.scala 12:21]
  wire  _T_241; // @[Shift.scala 12:21]
  wire [1:0] _T_243; // @[Bitwise.scala 71:12]
  wire [6:0] _T_244; // @[Cat.scala 29:58]
  wire [6:0] _T_245; // @[Shift.scala 91:22]
  wire  _T_246; // @[Shift.scala 92:77]
  wire [5:0] _T_247; // @[Shift.scala 90:30]
  wire  _T_248; // @[Shift.scala 90:48]
  wire [5:0] _GEN_16; // @[Shift.scala 90:39]
  wire [5:0] _T_250; // @[Shift.scala 90:39]
  wire  _T_252; // @[Shift.scala 12:21]
  wire [6:0] _T_253; // @[Cat.scala 29:58]
  wire [6:0] _T_254; // @[Shift.scala 91:22]
  wire [6:0] _T_257; // @[Bitwise.scala 71:12]
  wire [6:0] smallerSig; // @[Shift.scala 39:10]
  wire [7:0] rawSumSig; // @[PositFMA.scala 119:34]
  wire  _T_258; // @[PositFMA.scala 120:42]
  wire  _T_259; // @[PositFMA.scala 120:46]
  wire  _T_260; // @[PositFMA.scala 120:79]
  wire  sumSign; // @[PositFMA.scala 120:63]
  wire [6:0] _T_262; // @[PositFMA.scala 121:50]
  wire [7:0] signSumSig; // @[Cat.scala 29:58]
  wire [6:0] _T_263; // @[PositFMA.scala 126:33]
  wire [6:0] _T_264; // @[PositFMA.scala 126:68]
  wire [6:0] sumXor; // @[PositFMA.scala 126:51]
  wire [3:0] _T_265; // @[LZD.scala 43:32]
  wire [1:0] _T_266; // @[LZD.scala 43:32]
  wire  _T_267; // @[LZD.scala 39:14]
  wire  _T_268; // @[LZD.scala 39:21]
  wire  _T_269; // @[LZD.scala 39:30]
  wire  _T_270; // @[LZD.scala 39:27]
  wire  _T_271; // @[LZD.scala 39:25]
  wire [1:0] _T_272; // @[Cat.scala 29:58]
  wire [1:0] _T_273; // @[LZD.scala 44:32]
  wire  _T_274; // @[LZD.scala 39:14]
  wire  _T_275; // @[LZD.scala 39:21]
  wire  _T_276; // @[LZD.scala 39:30]
  wire  _T_277; // @[LZD.scala 39:27]
  wire  _T_278; // @[LZD.scala 39:25]
  wire [1:0] _T_279; // @[Cat.scala 29:58]
  wire  _T_280; // @[Shift.scala 12:21]
  wire  _T_281; // @[Shift.scala 12:21]
  wire  _T_282; // @[LZD.scala 49:16]
  wire  _T_283; // @[LZD.scala 49:27]
  wire  _T_284; // @[LZD.scala 49:25]
  wire  _T_285; // @[LZD.scala 49:47]
  wire  _T_286; // @[LZD.scala 49:59]
  wire  _T_287; // @[LZD.scala 49:35]
  wire [2:0] _T_289; // @[Cat.scala 29:58]
  wire [2:0] _T_290; // @[LZD.scala 44:32]
  wire [1:0] _T_291; // @[LZD.scala 43:32]
  wire  _T_292; // @[LZD.scala 39:14]
  wire  _T_293; // @[LZD.scala 39:21]
  wire  _T_294; // @[LZD.scala 39:30]
  wire  _T_295; // @[LZD.scala 39:27]
  wire  _T_296; // @[LZD.scala 39:25]
  wire [1:0] _T_297; // @[Cat.scala 29:58]
  wire  _T_298; // @[LZD.scala 44:32]
  wire  _T_300; // @[Shift.scala 12:21]
  wire  _T_302; // @[LZD.scala 55:32]
  wire  _T_303; // @[LZD.scala 55:20]
  wire [1:0] _T_304; // @[Cat.scala 29:58]
  wire  _T_305; // @[Shift.scala 12:21]
  wire [1:0] _T_307; // @[LZD.scala 55:32]
  wire [1:0] _T_308; // @[LZD.scala 55:20]
  wire [2:0] sumLZD; // @[Cat.scala 29:58]
  wire [2:0] shiftValue; // @[PositFMA.scala 128:24]
  wire [5:0] _T_309; // @[PositFMA.scala 129:38]
  wire  _T_310; // @[Shift.scala 16:24]
  wire  _T_312; // @[Shift.scala 12:21]
  wire [1:0] _T_313; // @[Shift.scala 64:52]
  wire [5:0] _T_315; // @[Cat.scala 29:58]
  wire [5:0] _T_316; // @[Shift.scala 64:27]
  wire [1:0] _T_317; // @[Shift.scala 66:70]
  wire  _T_318; // @[Shift.scala 12:21]
  wire [3:0] _T_319; // @[Shift.scala 64:52]
  wire [5:0] _T_321; // @[Cat.scala 29:58]
  wire [5:0] _T_322; // @[Shift.scala 64:27]
  wire  _T_323; // @[Shift.scala 66:70]
  wire [4:0] _T_325; // @[Shift.scala 64:52]
  wire [5:0] _T_326; // @[Cat.scala 29:58]
  wire [5:0] _T_327; // @[Shift.scala 64:27]
  wire [5:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [3:0] _T_329; // @[PositFMA.scala 132:36]
  wire [3:0] _T_330; // @[PositFMA.scala 132:36]
  wire [3:0] _T_331; // @[Cat.scala 29:58]
  wire [3:0] _T_332; // @[PositFMA.scala 132:61]
  wire [3:0] _T_334; // @[PositFMA.scala 132:42]
  wire [3:0] sumScale; // @[PositFMA.scala 132:42]
  wire [1:0] sumFrac; // @[PositFMA.scala 133:41]
  wire [3:0] grsTmp; // @[PositFMA.scala 136:41]
  wire [1:0] _T_335; // @[PositFMA.scala 139:40]
  wire [1:0] _T_336; // @[PositFMA.scala 139:56]
  wire  _T_337; // @[PositFMA.scala 139:60]
  wire  underflow; // @[PositFMA.scala 146:32]
  wire  overflow; // @[PositFMA.scala 147:32]
  wire  _T_338; // @[PositFMA.scala 156:32]
  wire  decF_isZero; // @[PositFMA.scala 156:20]
  wire [3:0] _T_340; // @[Mux.scala 87:16]
  wire [3:0] _T_341; // @[Mux.scala 87:16]
  wire [2:0] _GEN_17; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  wire [2:0] decF_scale; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  wire  _T_343; // @[convert.scala 49:36]
  wire [2:0] _T_345; // @[convert.scala 50:36]
  wire [2:0] _T_346; // @[convert.scala 50:36]
  wire [2:0] _T_347; // @[convert.scala 50:28]
  wire  _T_348; // @[convert.scala 51:31]
  wire  _T_349; // @[convert.scala 53:34]
  wire [6:0] _T_352; // @[Cat.scala 29:58]
  wire [2:0] _T_353; // @[Shift.scala 39:17]
  wire  _T_354; // @[Shift.scala 39:24]
  wire [2:0] _T_356; // @[Shift.scala 90:30]
  wire [3:0] _T_357; // @[Shift.scala 90:48]
  wire  _T_358; // @[Shift.scala 90:57]
  wire [2:0] _GEN_18; // @[Shift.scala 90:39]
  wire [2:0] _T_359; // @[Shift.scala 90:39]
  wire  _T_360; // @[Shift.scala 12:21]
  wire  _T_361; // @[Shift.scala 12:21]
  wire [3:0] _T_363; // @[Bitwise.scala 71:12]
  wire [6:0] _T_364; // @[Cat.scala 29:58]
  wire [6:0] _T_365; // @[Shift.scala 91:22]
  wire [1:0] _T_366; // @[Shift.scala 92:77]
  wire [4:0] _T_367; // @[Shift.scala 90:30]
  wire [1:0] _T_368; // @[Shift.scala 90:48]
  wire  _T_369; // @[Shift.scala 90:57]
  wire [4:0] _GEN_19; // @[Shift.scala 90:39]
  wire [4:0] _T_370; // @[Shift.scala 90:39]
  wire  _T_371; // @[Shift.scala 12:21]
  wire  _T_372; // @[Shift.scala 12:21]
  wire [1:0] _T_374; // @[Bitwise.scala 71:12]
  wire [6:0] _T_375; // @[Cat.scala 29:58]
  wire [6:0] _T_376; // @[Shift.scala 91:22]
  wire  _T_377; // @[Shift.scala 92:77]
  wire [5:0] _T_378; // @[Shift.scala 90:30]
  wire  _T_379; // @[Shift.scala 90:48]
  wire [5:0] _GEN_20; // @[Shift.scala 90:39]
  wire [5:0] _T_381; // @[Shift.scala 90:39]
  wire  _T_383; // @[Shift.scala 12:21]
  wire [6:0] _T_384; // @[Cat.scala 29:58]
  wire [6:0] _T_385; // @[Shift.scala 91:22]
  wire [6:0] _T_388; // @[Bitwise.scala 71:12]
  wire [6:0] _T_389; // @[Shift.scala 39:10]
  wire  _T_390; // @[convert.scala 55:31]
  wire  _T_391; // @[convert.scala 56:31]
  wire  _T_392; // @[convert.scala 57:31]
  wire  _T_393; // @[convert.scala 58:31]
  wire [3:0] _T_394; // @[convert.scala 59:69]
  wire  _T_395; // @[convert.scala 59:81]
  wire  _T_396; // @[convert.scala 59:50]
  wire  _T_398; // @[convert.scala 60:81]
  wire  _T_399; // @[convert.scala 61:44]
  wire  _T_400; // @[convert.scala 61:52]
  wire  _T_401; // @[convert.scala 61:36]
  wire  _T_402; // @[convert.scala 62:63]
  wire  _T_403; // @[convert.scala 62:103]
  wire  _T_404; // @[convert.scala 62:60]
  wire [3:0] _GEN_21; // @[convert.scala 63:56]
  wire [3:0] _T_407; // @[convert.scala 63:56]
  wire [4:0] _T_408; // @[Cat.scala 29:58]
  reg  _T_412; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [4:0] _T_416; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 5'h1f : 5'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{4'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 5'h1f : 5'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{4'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[4]; // @[convert.scala 18:24]
  assign _T_14 = realA[3]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[3:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[2:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[2:1]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19 != 2'h0; // @[LZD.scala 39:14]
  assign _T_21 = _T_19[1]; // @[LZD.scala 39:21]
  assign _T_22 = _T_19[0]; // @[LZD.scala 39:30]
  assign _T_23 = ~ _T_22; // @[LZD.scala 39:27]
  assign _T_24 = _T_21 | _T_23; // @[LZD.scala 39:25]
  assign _T_25 = {_T_20,_T_24}; // @[Cat.scala 29:58]
  assign _T_26 = _T_18[0:0]; // @[LZD.scala 44:32]
  assign _T_28 = _T_25[1]; // @[Shift.scala 12:21]
  assign _T_30 = _T_25[0:0]; // @[LZD.scala 55:32]
  assign _T_31 = _T_28 ? _T_30 : _T_26; // @[LZD.scala 55:20]
  assign _T_32 = {_T_28,_T_31}; // @[Cat.scala 29:58]
  assign _T_33 = ~ _T_32; // @[convert.scala 21:22]
  assign _T_34 = realA[1:0]; // @[convert.scala 22:36]
  assign _T_35 = _T_33 < 2'h2; // @[Shift.scala 16:24]
  assign _T_36 = _T_33[0]; // @[Shift.scala 17:37]
  assign _T_38 = _T_34[0:0]; // @[Shift.scala 64:52]
  assign _T_39 = {_T_38,1'h0}; // @[Cat.scala 29:58]
  assign _T_40 = _T_36 ? _T_39 : _T_34; // @[Shift.scala 64:27]
  assign decA_fraction = _T_35 ? _T_40 : 2'h0; // @[Shift.scala 16:10]
  assign _T_44 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_46 = _T_15 ? _T_33 : _T_32; // @[convert.scala 25:42]
  assign _T_47 = {_T_44,_T_46}; // @[Cat.scala 29:58]
  assign _T_49 = realA[3:0]; // @[convert.scala 29:56]
  assign _T_50 = _T_49 != 4'h0; // @[convert.scala 29:60]
  assign _T_51 = ~ _T_50; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_51; // @[convert.scala 29:39]
  assign _T_54 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_54 & _T_51; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_47); // @[convert.scala 32:24]
  assign _T_63 = io_B[4]; // @[convert.scala 18:24]
  assign _T_64 = io_B[3]; // @[convert.scala 18:40]
  assign _T_65 = _T_63 ^ _T_64; // @[convert.scala 18:36]
  assign _T_66 = io_B[3:1]; // @[convert.scala 19:24]
  assign _T_67 = io_B[2:0]; // @[convert.scala 19:43]
  assign _T_68 = _T_66 ^ _T_67; // @[convert.scala 19:39]
  assign _T_69 = _T_68[2:1]; // @[LZD.scala 43:32]
  assign _T_70 = _T_69 != 2'h0; // @[LZD.scala 39:14]
  assign _T_71 = _T_69[1]; // @[LZD.scala 39:21]
  assign _T_72 = _T_69[0]; // @[LZD.scala 39:30]
  assign _T_73 = ~ _T_72; // @[LZD.scala 39:27]
  assign _T_74 = _T_71 | _T_73; // @[LZD.scala 39:25]
  assign _T_75 = {_T_70,_T_74}; // @[Cat.scala 29:58]
  assign _T_76 = _T_68[0:0]; // @[LZD.scala 44:32]
  assign _T_78 = _T_75[1]; // @[Shift.scala 12:21]
  assign _T_80 = _T_75[0:0]; // @[LZD.scala 55:32]
  assign _T_81 = _T_78 ? _T_80 : _T_76; // @[LZD.scala 55:20]
  assign _T_82 = {_T_78,_T_81}; // @[Cat.scala 29:58]
  assign _T_83 = ~ _T_82; // @[convert.scala 21:22]
  assign _T_84 = io_B[1:0]; // @[convert.scala 22:36]
  assign _T_85 = _T_83 < 2'h2; // @[Shift.scala 16:24]
  assign _T_86 = _T_83[0]; // @[Shift.scala 17:37]
  assign _T_88 = _T_84[0:0]; // @[Shift.scala 64:52]
  assign _T_89 = {_T_88,1'h0}; // @[Cat.scala 29:58]
  assign _T_90 = _T_86 ? _T_89 : _T_84; // @[Shift.scala 64:27]
  assign decB_fraction = _T_85 ? _T_90 : 2'h0; // @[Shift.scala 16:10]
  assign _T_94 = _T_65 == 1'h0; // @[convert.scala 25:26]
  assign _T_96 = _T_65 ? _T_83 : _T_82; // @[convert.scala 25:42]
  assign _T_97 = {_T_94,_T_96}; // @[Cat.scala 29:58]
  assign _T_99 = io_B[3:0]; // @[convert.scala 29:56]
  assign _T_100 = _T_99 != 4'h0; // @[convert.scala 29:60]
  assign _T_101 = ~ _T_100; // @[convert.scala 29:41]
  assign decB_isNaR = _T_63 & _T_101; // @[convert.scala 29:39]
  assign _T_104 = _T_63 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_104 & _T_101; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_97); // @[convert.scala 32:24]
  assign _T_113 = realC[4]; // @[convert.scala 18:24]
  assign _T_114 = realC[3]; // @[convert.scala 18:40]
  assign _T_115 = _T_113 ^ _T_114; // @[convert.scala 18:36]
  assign _T_116 = realC[3:1]; // @[convert.scala 19:24]
  assign _T_117 = realC[2:0]; // @[convert.scala 19:43]
  assign _T_118 = _T_116 ^ _T_117; // @[convert.scala 19:39]
  assign _T_119 = _T_118[2:1]; // @[LZD.scala 43:32]
  assign _T_120 = _T_119 != 2'h0; // @[LZD.scala 39:14]
  assign _T_121 = _T_119[1]; // @[LZD.scala 39:21]
  assign _T_122 = _T_119[0]; // @[LZD.scala 39:30]
  assign _T_123 = ~ _T_122; // @[LZD.scala 39:27]
  assign _T_124 = _T_121 | _T_123; // @[LZD.scala 39:25]
  assign _T_125 = {_T_120,_T_124}; // @[Cat.scala 29:58]
  assign _T_126 = _T_118[0:0]; // @[LZD.scala 44:32]
  assign _T_128 = _T_125[1]; // @[Shift.scala 12:21]
  assign _T_130 = _T_125[0:0]; // @[LZD.scala 55:32]
  assign _T_131 = _T_128 ? _T_130 : _T_126; // @[LZD.scala 55:20]
  assign _T_132 = {_T_128,_T_131}; // @[Cat.scala 29:58]
  assign _T_133 = ~ _T_132; // @[convert.scala 21:22]
  assign _T_134 = realC[1:0]; // @[convert.scala 22:36]
  assign _T_135 = _T_133 < 2'h2; // @[Shift.scala 16:24]
  assign _T_136 = _T_133[0]; // @[Shift.scala 17:37]
  assign _T_138 = _T_134[0:0]; // @[Shift.scala 64:52]
  assign _T_139 = {_T_138,1'h0}; // @[Cat.scala 29:58]
  assign _T_144 = _T_115 == 1'h0; // @[convert.scala 25:26]
  assign _T_146 = _T_115 ? _T_133 : _T_132; // @[convert.scala 25:42]
  assign _T_147 = {_T_144,_T_146}; // @[Cat.scala 29:58]
  assign _T_149 = realC[3:0]; // @[convert.scala 29:56]
  assign _T_150 = _T_149 != 4'h0; // @[convert.scala 29:60]
  assign _T_151 = ~ _T_150; // @[convert.scala 29:41]
  assign decC_isNaR = _T_113 & _T_151; // @[convert.scala 29:39]
  assign _T_154 = _T_113 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_154 & _T_151; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_147); // @[convert.scala 32:24]
  assign _T_162 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_162 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_163 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_164 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_165 = _T_163 & _T_164; // @[PositFMA.scala 59:45]
  assign _T_167 = {_T_13,_T_165,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_167); // @[PositFMA.scala 59:76]
  assign _T_168 = ~ _T_63; // @[PositFMA.scala 60:34]
  assign _T_169 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_170 = _T_168 & _T_169; // @[PositFMA.scala 60:45]
  assign _T_172 = {_T_63,_T_170,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_172); // @[PositFMA.scala 60:76]
  assign _T_173 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 62:25]
  assign sigP = $unsigned(_T_173); // @[PositFMA.scala 62:33]
  assign head2 = sigP[7:6]; // @[PositFMA.scala 63:28]
  assign _T_174 = head2[1]; // @[PositFMA.scala 64:31]
  assign _T_175 = ~ _T_174; // @[PositFMA.scala 64:25]
  assign _T_176 = head2[0]; // @[PositFMA.scala 64:42]
  assign addTwo = _T_175 & _T_176; // @[PositFMA.scala 64:35]
  assign _T_177 = sigP[7]; // @[PositFMA.scala 66:23]
  assign _T_178 = sigP[5]; // @[PositFMA.scala 66:49]
  assign addOne = _T_177 ^ _T_178; // @[PositFMA.scala 66:43]
  assign _T_179 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_179)}; // @[PositFMA.scala 67:39]
  assign mulSign = sigP[7:7]; // @[PositFMA.scala 68:28]
  assign _T_180 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 70:30]
  assign _GEN_12 = {{1{expBias[2]}},expBias}; // @[PositFMA.scala 70:44]
  assign _T_182 = $signed(_T_180) + $signed(_GEN_12); // @[PositFMA.scala 70:44]
  assign mulScale = $signed(_T_182); // @[PositFMA.scala 70:44]
  assign _T_183 = sigP[5:0]; // @[PositFMA.scala 73:29]
  assign _T_184 = sigP[4:0]; // @[PositFMA.scala 74:29]
  assign _T_185 = {_T_184, 1'h0}; // @[PositFMA.scala 74:48]
  assign mulSigTmp = addOne ? _T_183 : _T_185; // @[PositFMA.scala 71:22]
  assign _T_187 = mulSigTmp[5:5]; // @[PositFMA.scala 78:39]
  assign _T_188 = _T_187 | addTwo; // @[PositFMA.scala 78:43]
  assign _T_189 = mulSigTmp[4:0]; // @[PositFMA.scala 79:39]
  assign mulSig = {mulSign,_T_188,_T_189}; // @[Cat.scala 29:58]
  assign _T_215 = ~ addSign_phase2; // @[PositFMA.scala 108:29]
  assign _T_216 = ~ addZero_phase2; // @[PositFMA.scala 108:47]
  assign _T_217 = _T_215 & _T_216; // @[PositFMA.scala 108:45]
  assign extAddSig = {addSign_phase2,_T_217,addFrac_phase2,3'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[2]}},addScale_phase2}; // @[PositFMA.scala 112:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 112:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[2]}},addScale_phase2}); // @[PositFMA.scala 113:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[2]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 114:26]
  assign _T_221 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 115:36]
  assign scaleDiff = $signed(_T_221); // @[PositFMA.scala 115:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 116:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 117:26]
  assign _T_222 = $unsigned(scaleDiff); // @[PositFMA.scala 118:69]
  assign _T_223 = _T_222 < 4'h7; // @[Shift.scala 39:24]
  assign _T_224 = _T_222[2:0]; // @[Shift.scala 40:44]
  assign _T_225 = smallerSigTmp[6:4]; // @[Shift.scala 90:30]
  assign _T_226 = smallerSigTmp[3:0]; // @[Shift.scala 90:48]
  assign _T_227 = _T_226 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{2'd0}, _T_227}; // @[Shift.scala 90:39]
  assign _T_228 = _T_225 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_229 = _T_224[2]; // @[Shift.scala 12:21]
  assign _T_230 = smallerSigTmp[6]; // @[Shift.scala 12:21]
  assign _T_232 = _T_230 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_233 = {_T_232,_T_228}; // @[Cat.scala 29:58]
  assign _T_234 = _T_229 ? _T_233 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_235 = _T_224[1:0]; // @[Shift.scala 92:77]
  assign _T_236 = _T_234[6:2]; // @[Shift.scala 90:30]
  assign _T_237 = _T_234[1:0]; // @[Shift.scala 90:48]
  assign _T_238 = _T_237 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{4'd0}, _T_238}; // @[Shift.scala 90:39]
  assign _T_239 = _T_236 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_240 = _T_235[1]; // @[Shift.scala 12:21]
  assign _T_241 = _T_234[6]; // @[Shift.scala 12:21]
  assign _T_243 = _T_241 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_244 = {_T_243,_T_239}; // @[Cat.scala 29:58]
  assign _T_245 = _T_240 ? _T_244 : _T_234; // @[Shift.scala 91:22]
  assign _T_246 = _T_235[0:0]; // @[Shift.scala 92:77]
  assign _T_247 = _T_245[6:1]; // @[Shift.scala 90:30]
  assign _T_248 = _T_245[0:0]; // @[Shift.scala 90:48]
  assign _GEN_16 = {{5'd0}, _T_248}; // @[Shift.scala 90:39]
  assign _T_250 = _T_247 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_252 = _T_245[6]; // @[Shift.scala 12:21]
  assign _T_253 = {_T_252,_T_250}; // @[Cat.scala 29:58]
  assign _T_254 = _T_246 ? _T_253 : _T_245; // @[Shift.scala 91:22]
  assign _T_257 = _T_230 ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_223 ? _T_254 : _T_257; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 119:34]
  assign _T_258 = mulSig_phase2[6:6]; // @[PositFMA.scala 120:42]
  assign _T_259 = _T_258 ^ addSign_phase2; // @[PositFMA.scala 120:46]
  assign _T_260 = rawSumSig[7:7]; // @[PositFMA.scala 120:79]
  assign sumSign = _T_259 ^ _T_260; // @[PositFMA.scala 120:63]
  assign _T_262 = greaterSig + smallerSig; // @[PositFMA.scala 121:50]
  assign signSumSig = {sumSign,_T_262}; // @[Cat.scala 29:58]
  assign _T_263 = signSumSig[7:1]; // @[PositFMA.scala 126:33]
  assign _T_264 = signSumSig[6:0]; // @[PositFMA.scala 126:68]
  assign sumXor = _T_263 ^ _T_264; // @[PositFMA.scala 126:51]
  assign _T_265 = sumXor[6:3]; // @[LZD.scala 43:32]
  assign _T_266 = _T_265[3:2]; // @[LZD.scala 43:32]
  assign _T_267 = _T_266 != 2'h0; // @[LZD.scala 39:14]
  assign _T_268 = _T_266[1]; // @[LZD.scala 39:21]
  assign _T_269 = _T_266[0]; // @[LZD.scala 39:30]
  assign _T_270 = ~ _T_269; // @[LZD.scala 39:27]
  assign _T_271 = _T_268 | _T_270; // @[LZD.scala 39:25]
  assign _T_272 = {_T_267,_T_271}; // @[Cat.scala 29:58]
  assign _T_273 = _T_265[1:0]; // @[LZD.scala 44:32]
  assign _T_274 = _T_273 != 2'h0; // @[LZD.scala 39:14]
  assign _T_275 = _T_273[1]; // @[LZD.scala 39:21]
  assign _T_276 = _T_273[0]; // @[LZD.scala 39:30]
  assign _T_277 = ~ _T_276; // @[LZD.scala 39:27]
  assign _T_278 = _T_275 | _T_277; // @[LZD.scala 39:25]
  assign _T_279 = {_T_274,_T_278}; // @[Cat.scala 29:58]
  assign _T_280 = _T_272[1]; // @[Shift.scala 12:21]
  assign _T_281 = _T_279[1]; // @[Shift.scala 12:21]
  assign _T_282 = _T_280 | _T_281; // @[LZD.scala 49:16]
  assign _T_283 = ~ _T_281; // @[LZD.scala 49:27]
  assign _T_284 = _T_280 | _T_283; // @[LZD.scala 49:25]
  assign _T_285 = _T_272[0:0]; // @[LZD.scala 49:47]
  assign _T_286 = _T_279[0:0]; // @[LZD.scala 49:59]
  assign _T_287 = _T_280 ? _T_285 : _T_286; // @[LZD.scala 49:35]
  assign _T_289 = {_T_282,_T_284,_T_287}; // @[Cat.scala 29:58]
  assign _T_290 = sumXor[2:0]; // @[LZD.scala 44:32]
  assign _T_291 = _T_290[2:1]; // @[LZD.scala 43:32]
  assign _T_292 = _T_291 != 2'h0; // @[LZD.scala 39:14]
  assign _T_293 = _T_291[1]; // @[LZD.scala 39:21]
  assign _T_294 = _T_291[0]; // @[LZD.scala 39:30]
  assign _T_295 = ~ _T_294; // @[LZD.scala 39:27]
  assign _T_296 = _T_293 | _T_295; // @[LZD.scala 39:25]
  assign _T_297 = {_T_292,_T_296}; // @[Cat.scala 29:58]
  assign _T_298 = _T_290[0:0]; // @[LZD.scala 44:32]
  assign _T_300 = _T_297[1]; // @[Shift.scala 12:21]
  assign _T_302 = _T_297[0:0]; // @[LZD.scala 55:32]
  assign _T_303 = _T_300 ? _T_302 : _T_298; // @[LZD.scala 55:20]
  assign _T_304 = {_T_300,_T_303}; // @[Cat.scala 29:58]
  assign _T_305 = _T_289[2]; // @[Shift.scala 12:21]
  assign _T_307 = _T_289[1:0]; // @[LZD.scala 55:32]
  assign _T_308 = _T_305 ? _T_307 : _T_304; // @[LZD.scala 55:20]
  assign sumLZD = {_T_305,_T_308}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 128:24]
  assign _T_309 = signSumSig[5:0]; // @[PositFMA.scala 129:38]
  assign _T_310 = shiftValue < 3'h6; // @[Shift.scala 16:24]
  assign _T_312 = shiftValue[2]; // @[Shift.scala 12:21]
  assign _T_313 = _T_309[1:0]; // @[Shift.scala 64:52]
  assign _T_315 = {_T_313,4'h0}; // @[Cat.scala 29:58]
  assign _T_316 = _T_312 ? _T_315 : _T_309; // @[Shift.scala 64:27]
  assign _T_317 = shiftValue[1:0]; // @[Shift.scala 66:70]
  assign _T_318 = _T_317[1]; // @[Shift.scala 12:21]
  assign _T_319 = _T_316[3:0]; // @[Shift.scala 64:52]
  assign _T_321 = {_T_319,2'h0}; // @[Cat.scala 29:58]
  assign _T_322 = _T_318 ? _T_321 : _T_316; // @[Shift.scala 64:27]
  assign _T_323 = _T_317[0:0]; // @[Shift.scala 66:70]
  assign _T_325 = _T_322[4:0]; // @[Shift.scala 64:52]
  assign _T_326 = {_T_325,1'h0}; // @[Cat.scala 29:58]
  assign _T_327 = _T_323 ? _T_326 : _T_322; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_310 ? _T_327 : 6'h0; // @[Shift.scala 16:10]
  assign _T_329 = $signed(greaterScale) + $signed(4'sh2); // @[PositFMA.scala 132:36]
  assign _T_330 = $signed(_T_329); // @[PositFMA.scala 132:36]
  assign _T_331 = {1'h1,_T_305,_T_308}; // @[Cat.scala 29:58]
  assign _T_332 = $signed(_T_331); // @[PositFMA.scala 132:61]
  assign _T_334 = $signed(_T_330) + $signed(_T_332); // @[PositFMA.scala 132:42]
  assign sumScale = $signed(_T_334); // @[PositFMA.scala 132:42]
  assign sumFrac = normalFracTmp[5:4]; // @[PositFMA.scala 133:41]
  assign grsTmp = normalFracTmp[3:0]; // @[PositFMA.scala 136:41]
  assign _T_335 = grsTmp[3:2]; // @[PositFMA.scala 139:40]
  assign _T_336 = grsTmp[1:0]; // @[PositFMA.scala 139:56]
  assign _T_337 = _T_336 != 2'h0; // @[PositFMA.scala 139:60]
  assign underflow = $signed(sumScale) < $signed(-4'sh4); // @[PositFMA.scala 146:32]
  assign overflow = $signed(sumScale) > $signed(4'sh3); // @[PositFMA.scala 147:32]
  assign _T_338 = signSumSig != 8'h0; // @[PositFMA.scala 156:32]
  assign decF_isZero = ~ _T_338; // @[PositFMA.scala 156:20]
  assign _T_340 = underflow ? $signed(-4'sh4) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_341 = overflow ? $signed(4'sh3) : $signed(_T_340); // @[Mux.scala 87:16]
  assign _GEN_17 = _T_341[2:0]; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  assign decF_scale = $signed(_GEN_17); // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  assign _T_343 = decF_scale[2:2]; // @[convert.scala 49:36]
  assign _T_345 = ~ decF_scale; // @[convert.scala 50:36]
  assign _T_346 = $signed(_T_345); // @[convert.scala 50:36]
  assign _T_347 = _T_343 ? $signed(_T_346) : $signed(decF_scale); // @[convert.scala 50:28]
  assign _T_348 = _T_343 ^ sumSign; // @[convert.scala 51:31]
  assign _T_349 = ~ _T_348; // @[convert.scala 53:34]
  assign _T_352 = {_T_349,_T_348,sumFrac,_T_335,_T_337}; // @[Cat.scala 29:58]
  assign _T_353 = $unsigned(_T_347); // @[Shift.scala 39:17]
  assign _T_354 = _T_353 < 3'h7; // @[Shift.scala 39:24]
  assign _T_356 = _T_352[6:4]; // @[Shift.scala 90:30]
  assign _T_357 = _T_352[3:0]; // @[Shift.scala 90:48]
  assign _T_358 = _T_357 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_18 = {{2'd0}, _T_358}; // @[Shift.scala 90:39]
  assign _T_359 = _T_356 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_360 = _T_353[2]; // @[Shift.scala 12:21]
  assign _T_361 = _T_352[6]; // @[Shift.scala 12:21]
  assign _T_363 = _T_361 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_364 = {_T_363,_T_359}; // @[Cat.scala 29:58]
  assign _T_365 = _T_360 ? _T_364 : _T_352; // @[Shift.scala 91:22]
  assign _T_366 = _T_353[1:0]; // @[Shift.scala 92:77]
  assign _T_367 = _T_365[6:2]; // @[Shift.scala 90:30]
  assign _T_368 = _T_365[1:0]; // @[Shift.scala 90:48]
  assign _T_369 = _T_368 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_19 = {{4'd0}, _T_369}; // @[Shift.scala 90:39]
  assign _T_370 = _T_367 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_371 = _T_366[1]; // @[Shift.scala 12:21]
  assign _T_372 = _T_365[6]; // @[Shift.scala 12:21]
  assign _T_374 = _T_372 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_375 = {_T_374,_T_370}; // @[Cat.scala 29:58]
  assign _T_376 = _T_371 ? _T_375 : _T_365; // @[Shift.scala 91:22]
  assign _T_377 = _T_366[0:0]; // @[Shift.scala 92:77]
  assign _T_378 = _T_376[6:1]; // @[Shift.scala 90:30]
  assign _T_379 = _T_376[0:0]; // @[Shift.scala 90:48]
  assign _GEN_20 = {{5'd0}, _T_379}; // @[Shift.scala 90:39]
  assign _T_381 = _T_378 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_383 = _T_376[6]; // @[Shift.scala 12:21]
  assign _T_384 = {_T_383,_T_381}; // @[Cat.scala 29:58]
  assign _T_385 = _T_377 ? _T_384 : _T_376; // @[Shift.scala 91:22]
  assign _T_388 = _T_361 ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign _T_389 = _T_354 ? _T_385 : _T_388; // @[Shift.scala 39:10]
  assign _T_390 = _T_389[3]; // @[convert.scala 55:31]
  assign _T_391 = _T_389[2]; // @[convert.scala 56:31]
  assign _T_392 = _T_389[1]; // @[convert.scala 57:31]
  assign _T_393 = _T_389[0]; // @[convert.scala 58:31]
  assign _T_394 = _T_389[6:3]; // @[convert.scala 59:69]
  assign _T_395 = _T_394 != 4'h0; // @[convert.scala 59:81]
  assign _T_396 = ~ _T_395; // @[convert.scala 59:50]
  assign _T_398 = _T_394 == 4'hf; // @[convert.scala 60:81]
  assign _T_399 = _T_390 | _T_392; // @[convert.scala 61:44]
  assign _T_400 = _T_399 | _T_393; // @[convert.scala 61:52]
  assign _T_401 = _T_391 & _T_400; // @[convert.scala 61:36]
  assign _T_402 = ~ _T_398; // @[convert.scala 62:63]
  assign _T_403 = _T_402 & _T_401; // @[convert.scala 62:103]
  assign _T_404 = _T_396 | _T_403; // @[convert.scala 62:60]
  assign _GEN_21 = {{3'd0}, _T_404}; // @[convert.scala 63:56]
  assign _T_407 = _T_394 + _GEN_21; // @[convert.scala 63:56]
  assign _T_408 = {sumSign,_T_407}; // @[Cat.scala 29:58]
  assign io_F = _T_416; // @[PositFMA.scala 176:15]
  assign io_outValid = _T_412; // @[PositFMA.scala 175:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulSig_phase2 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_412 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_416 = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      if (_T_135) begin
        if (_T_136) begin
          addFrac_phase2 <= _T_139;
        end else begin
          addFrac_phase2 <= _T_134;
        end
      end else begin
        addFrac_phase2 <= 2'h0;
      end
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_113;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_412 <= 1'h0;
    end else begin
      _T_412 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_416 <= 5'h10;
      end else begin
        if (decF_isZero) begin
          _T_416 <= 5'h0;
        end else begin
          _T_416 <= _T_408;
        end
      end
    end
  end
endmodule
