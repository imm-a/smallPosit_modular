module PositDivSqrter6_0(
  input        clock,
  input        reset,
  output       io_inReady,
  input        io_inValid,
  input        io_sqrtOp,
  input  [5:0] io_A,
  input  [5:0] io_B,
  output       io_diviValid,
  output       io_sqrtValid,
  output       io_invalidExc,
  output [5:0] io_Q
);
  reg [3:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [4:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg [2:0] fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [9:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [9:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [3:0] _T_4; // @[convert.scala 19:24]
  wire [3:0] _T_5; // @[convert.scala 19:43]
  wire [3:0] _T_6; // @[convert.scala 19:39]
  wire [1:0] _T_7; // @[LZD.scala 43:32]
  wire  _T_8; // @[LZD.scala 39:14]
  wire  _T_9; // @[LZD.scala 39:21]
  wire  _T_10; // @[LZD.scala 39:30]
  wire  _T_11; // @[LZD.scala 39:27]
  wire  _T_12; // @[LZD.scala 39:25]
  wire [1:0] _T_13; // @[Cat.scala 29:58]
  wire [1:0] _T_14; // @[LZD.scala 44:32]
  wire  _T_15; // @[LZD.scala 39:14]
  wire  _T_16; // @[LZD.scala 39:21]
  wire  _T_17; // @[LZD.scala 39:30]
  wire  _T_18; // @[LZD.scala 39:27]
  wire  _T_19; // @[LZD.scala 39:25]
  wire [1:0] _T_20; // @[Cat.scala 29:58]
  wire  _T_21; // @[Shift.scala 12:21]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[LZD.scala 49:16]
  wire  _T_24; // @[LZD.scala 49:27]
  wire  _T_25; // @[LZD.scala 49:25]
  wire  _T_26; // @[LZD.scala 49:47]
  wire  _T_27; // @[LZD.scala 49:59]
  wire  _T_28; // @[LZD.scala 49:35]
  wire [2:0] _T_30; // @[Cat.scala 29:58]
  wire [2:0] _T_31; // @[convert.scala 21:22]
  wire [2:0] _T_32; // @[convert.scala 22:36]
  wire  _T_33; // @[Shift.scala 16:24]
  wire [1:0] _T_34; // @[Shift.scala 17:37]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[Shift.scala 64:52]
  wire [2:0] _T_38; // @[Cat.scala 29:58]
  wire [2:0] _T_39; // @[Shift.scala 64:27]
  wire  _T_40; // @[Shift.scala 66:70]
  wire [1:0] _T_42; // @[Shift.scala 64:52]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire [2:0] _T_44; // @[Shift.scala 64:27]
  wire [2:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_48; // @[convert.scala 25:26]
  wire [2:0] _T_50; // @[convert.scala 25:42]
  wire [3:0] _T_51; // @[Cat.scala 29:58]
  wire [4:0] _T_53; // @[convert.scala 29:56]
  wire  _T_54; // @[convert.scala 29:60]
  wire  _T_55; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_58; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [3:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_67; // @[convert.scala 18:24]
  wire  _T_68; // @[convert.scala 18:40]
  wire  _T_69; // @[convert.scala 18:36]
  wire [3:0] _T_70; // @[convert.scala 19:24]
  wire [3:0] _T_71; // @[convert.scala 19:43]
  wire [3:0] _T_72; // @[convert.scala 19:39]
  wire [1:0] _T_73; // @[LZD.scala 43:32]
  wire  _T_74; // @[LZD.scala 39:14]
  wire  _T_75; // @[LZD.scala 39:21]
  wire  _T_76; // @[LZD.scala 39:30]
  wire  _T_77; // @[LZD.scala 39:27]
  wire  _T_78; // @[LZD.scala 39:25]
  wire [1:0] _T_79; // @[Cat.scala 29:58]
  wire [1:0] _T_80; // @[LZD.scala 44:32]
  wire  _T_81; // @[LZD.scala 39:14]
  wire  _T_82; // @[LZD.scala 39:21]
  wire  _T_83; // @[LZD.scala 39:30]
  wire  _T_84; // @[LZD.scala 39:27]
  wire  _T_85; // @[LZD.scala 39:25]
  wire [1:0] _T_86; // @[Cat.scala 29:58]
  wire  _T_87; // @[Shift.scala 12:21]
  wire  _T_88; // @[Shift.scala 12:21]
  wire  _T_89; // @[LZD.scala 49:16]
  wire  _T_90; // @[LZD.scala 49:27]
  wire  _T_91; // @[LZD.scala 49:25]
  wire  _T_92; // @[LZD.scala 49:47]
  wire  _T_93; // @[LZD.scala 49:59]
  wire  _T_94; // @[LZD.scala 49:35]
  wire [2:0] _T_96; // @[Cat.scala 29:58]
  wire [2:0] _T_97; // @[convert.scala 21:22]
  wire [2:0] _T_98; // @[convert.scala 22:36]
  wire  _T_99; // @[Shift.scala 16:24]
  wire [1:0] _T_100; // @[Shift.scala 17:37]
  wire  _T_101; // @[Shift.scala 12:21]
  wire  _T_102; // @[Shift.scala 64:52]
  wire [2:0] _T_104; // @[Cat.scala 29:58]
  wire [2:0] _T_105; // @[Shift.scala 64:27]
  wire  _T_106; // @[Shift.scala 66:70]
  wire [1:0] _T_108; // @[Shift.scala 64:52]
  wire [2:0] _T_109; // @[Cat.scala 29:58]
  wire [2:0] _T_110; // @[Shift.scala 64:27]
  wire [2:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_114; // @[convert.scala 25:26]
  wire [2:0] _T_116; // @[convert.scala 25:42]
  wire [3:0] _T_117; // @[Cat.scala 29:58]
  wire [4:0] _T_119; // @[convert.scala 29:56]
  wire  _T_120; // @[convert.scala 29:60]
  wire  _T_121; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_124; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [3:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_133; // @[Bitwise.scala 71:12]
  wire  _T_134; // @[PositDivisionSqrt.scala 80:40]
  wire [9:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_137; // @[PositDivisionSqrt.scala 82:31]
  wire [9:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_140; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_141; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_142; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_143; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_144; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_145; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_146; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_147; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_148; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_149; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [4:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_152; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_153; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_154; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_155; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_156; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_157; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_158; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_159; // @[PositDivisionSqrt.scala 117:30]
  wire [3:0] _T_161; // @[PositDivisionSqrt.scala 119:26]
  wire [3:0] _T_162; // @[PositDivisionSqrt.scala 118:20]
  wire [3:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [3:0] _T_163; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_165; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_166; // @[PositDivisionSqrt.scala 123:27]
  wire [3:0] _T_168; // @[PositDivisionSqrt.scala 123:52]
  wire [3:0] _T_169; // @[PositDivisionSqrt.scala 123:20]
  wire [3:0] _T_170; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_172; // @[PositDivisionSqrt.scala 124:27]
  wire [3:0] _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _T_174; // @[PositDivisionSqrt.scala 123:64]
  wire [2:0] _T_175; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_177; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_178; // @[PositDivisionSqrt.scala 137:28]
  wire [15:0] _T_179; // @[PositDivisionSqrt.scala 146:22]
  wire [13:0] _T_180; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_181; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_182; // @[PositDivisionSqrt.scala 148:23]
  wire [9:0] _T_183; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_184; // @[PositDivisionSqrt.scala 149:23]
  wire [10:0] _T_185; // @[PositDivisionSqrt.scala 149:46]
  wire [9:0] _T_186; // @[PositDivisionSqrt.scala 149:56]
  wire [9:0] _T_187; // @[PositDivisionSqrt.scala 149:16]
  wire [9:0] _T_188; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_189; // @[PositDivisionSqrt.scala 150:17]
  wire [9:0] _T_190; // @[PositDivisionSqrt.scala 150:16]
  wire [9:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_192; // @[PositDivisionSqrt.scala 152:29]
  wire [9:0] _T_193; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_194; // @[PositDivisionSqrt.scala 153:29]
  wire [6:0] _T_195; // @[PositDivisionSqrt.scala 153:22]
  wire [9:0] _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  wire [9:0] _T_196; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_198; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_199; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_200; // @[PositDivisionSqrt.scala 154:57]
  wire [9:0] _T_203; // @[Cat.scala 29:58]
  wire [9:0] _T_204; // @[PositDivisionSqrt.scala 154:22]
  wire [9:0] _T_205; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_207; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_208; // @[PositDivisionSqrt.scala 156:83]
  wire [5:0] _T_210; // @[Bitwise.scala 71:12]
  wire [8:0] bitMask; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  wire [8:0] _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  wire [8:0] _T_211; // @[PositDivisionSqrt.scala 156:53]
  wire [9:0] _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  wire [9:0] _T_212; // @[PositDivisionSqrt.scala 155:51]
  wire [7:0] _T_213; // @[PositDivisionSqrt.scala 157:53]
  wire [9:0] _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  wire [9:0] _T_214; // @[PositDivisionSqrt.scala 156:89]
  wire [9:0] _T_215; // @[PositDivisionSqrt.scala 155:22]
  wire [9:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_217; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_218; // @[PositDivisionSqrt.scala 162:40]
  wire [9:0] _T_221; // @[PositDivisionSqrt.scala 163:97]
  wire [9:0] _T_223; // @[PositDivisionSqrt.scala 164:97]
  wire [9:0] _T_224; // @[PositDivisionSqrt.scala 161:92]
  wire [10:0] _T_229; // @[PositDivisionSqrt.scala 168:98]
  wire [9:0] _T_230; // @[PositDivisionSqrt.scala 168:108]
  wire [9:0] _T_232; // @[PositDivisionSqrt.scala 168:112]
  wire [9:0] _T_236; // @[PositDivisionSqrt.scala 169:112]
  wire [9:0] _T_237; // @[PositDivisionSqrt.scala 166:26]
  wire [9:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_238; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_239; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_241; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_242; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_243; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_244; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_245; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_247; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_248; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_249; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_250; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_251; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_254; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_255; // @[PositDivisionSqrt.scala 187:28]
  wire [9:0] _T_258; // @[PositDivisionSqrt.scala 188:47]
  wire [9:0] _T_259; // @[PositDivisionSqrt.scala 188:18]
  wire [7:0] _T_261; // @[PositDivisionSqrt.scala 189:18]
  wire [9:0] _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  wire [9:0] _T_262; // @[PositDivisionSqrt.scala 188:78]
  wire [9:0] _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  wire [9:0] _T_264; // @[PositDivisionSqrt.scala 190:47]
  wire [9:0] _T_265; // @[PositDivisionSqrt.scala 190:18]
  wire [9:0] _T_266; // @[PositDivisionSqrt.scala 189:78]
  wire [1:0] _T_268; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [9:0] _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  wire [9:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire [2:0] _T_271; // @[PositDivisionSqrt.scala 200:97]
  wire [2:0] _T_272; // @[PositDivisionSqrt.scala 201:97]
  wire [2:0] realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_273; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_274; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_275; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  _T_277; // @[PositDivisionSqrt.scala 206:56]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_278; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_279; // @[Cat.scala 29:58]
  wire [2:0] _T_280; // @[PositDivisionSqrt.scala 209:63]
  wire [4:0] _GEN_18; // @[PositDivisionSqrt.scala 209:31]
  wire [4:0] _T_282; // @[PositDivisionSqrt.scala 209:31]
  wire [4:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [4:0] _T_284; // @[Mux.scala 87:16]
  wire [4:0] _T_285; // @[Mux.scala 87:16]
  wire [2:0] _T_286; // @[PositDivisionSqrt.scala 224:48]
  wire [2:0] _T_287; // @[PositDivisionSqrt.scala 224:64]
  wire [2:0] decQ_grs; // @[PositDivisionSqrt.scala 224:23]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [3:0] _GEN_19; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [3:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire  _T_294; // @[convert.scala 49:36]
  wire [3:0] _T_296; // @[convert.scala 50:36]
  wire [3:0] _T_297; // @[convert.scala 50:36]
  wire [3:0] _T_298; // @[convert.scala 50:28]
  wire  _T_299; // @[convert.scala 51:31]
  wire  _T_300; // @[convert.scala 53:34]
  wire [7:0] _T_303; // @[Cat.scala 29:58]
  wire [3:0] _T_304; // @[Shift.scala 39:17]
  wire  _T_305; // @[Shift.scala 39:24]
  wire [2:0] _T_306; // @[Shift.scala 40:44]
  wire [3:0] _T_307; // @[Shift.scala 90:30]
  wire [3:0] _T_308; // @[Shift.scala 90:48]
  wire  _T_309; // @[Shift.scala 90:57]
  wire [3:0] _GEN_20; // @[Shift.scala 90:39]
  wire [3:0] _T_310; // @[Shift.scala 90:39]
  wire  _T_311; // @[Shift.scala 12:21]
  wire  _T_312; // @[Shift.scala 12:21]
  wire [3:0] _T_314; // @[Bitwise.scala 71:12]
  wire [7:0] _T_315; // @[Cat.scala 29:58]
  wire [7:0] _T_316; // @[Shift.scala 91:22]
  wire [1:0] _T_317; // @[Shift.scala 92:77]
  wire [5:0] _T_318; // @[Shift.scala 90:30]
  wire [1:0] _T_319; // @[Shift.scala 90:48]
  wire  _T_320; // @[Shift.scala 90:57]
  wire [5:0] _GEN_21; // @[Shift.scala 90:39]
  wire [5:0] _T_321; // @[Shift.scala 90:39]
  wire  _T_322; // @[Shift.scala 12:21]
  wire  _T_323; // @[Shift.scala 12:21]
  wire [1:0] _T_325; // @[Bitwise.scala 71:12]
  wire [7:0] _T_326; // @[Cat.scala 29:58]
  wire [7:0] _T_327; // @[Shift.scala 91:22]
  wire  _T_328; // @[Shift.scala 92:77]
  wire [6:0] _T_329; // @[Shift.scala 90:30]
  wire  _T_330; // @[Shift.scala 90:48]
  wire [6:0] _GEN_22; // @[Shift.scala 90:39]
  wire [6:0] _T_332; // @[Shift.scala 90:39]
  wire  _T_334; // @[Shift.scala 12:21]
  wire [7:0] _T_335; // @[Cat.scala 29:58]
  wire [7:0] _T_336; // @[Shift.scala 91:22]
  wire [7:0] _T_339; // @[Bitwise.scala 71:12]
  wire [7:0] _T_340; // @[Shift.scala 39:10]
  wire  _T_341; // @[convert.scala 55:31]
  wire  _T_342; // @[convert.scala 56:31]
  wire  _T_343; // @[convert.scala 57:31]
  wire  _T_344; // @[convert.scala 58:31]
  wire [4:0] _T_345; // @[convert.scala 59:69]
  wire  _T_346; // @[convert.scala 59:81]
  wire  _T_347; // @[convert.scala 59:50]
  wire  _T_349; // @[convert.scala 60:81]
  wire  _T_350; // @[convert.scala 61:44]
  wire  _T_351; // @[convert.scala 61:52]
  wire  _T_352; // @[convert.scala 61:36]
  wire  _T_353; // @[convert.scala 62:63]
  wire  _T_354; // @[convert.scala 62:103]
  wire  _T_355; // @[convert.scala 62:60]
  wire [4:0] _GEN_23; // @[convert.scala 63:56]
  wire [4:0] _T_358; // @[convert.scala 63:56]
  wire [5:0] _T_359; // @[Cat.scala 29:58]
  wire [5:0] _T_361; // @[Mux.scala 87:16]
  assign _T_1 = io_A[5]; // @[convert.scala 18:24]
  assign _T_2 = io_A[4]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[4:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[3:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[3:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7 != 2'h0; // @[LZD.scala 39:14]
  assign _T_9 = _T_7[1]; // @[LZD.scala 39:21]
  assign _T_10 = _T_7[0]; // @[LZD.scala 39:30]
  assign _T_11 = ~ _T_10; // @[LZD.scala 39:27]
  assign _T_12 = _T_9 | _T_11; // @[LZD.scala 39:25]
  assign _T_13 = {_T_8,_T_12}; // @[Cat.scala 29:58]
  assign _T_14 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_15 = _T_14 != 2'h0; // @[LZD.scala 39:14]
  assign _T_16 = _T_14[1]; // @[LZD.scala 39:21]
  assign _T_17 = _T_14[0]; // @[LZD.scala 39:30]
  assign _T_18 = ~ _T_17; // @[LZD.scala 39:27]
  assign _T_19 = _T_16 | _T_18; // @[LZD.scala 39:25]
  assign _T_20 = {_T_15,_T_19}; // @[Cat.scala 29:58]
  assign _T_21 = _T_13[1]; // @[Shift.scala 12:21]
  assign _T_22 = _T_20[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21 | _T_22; // @[LZD.scala 49:16]
  assign _T_24 = ~ _T_22; // @[LZD.scala 49:27]
  assign _T_25 = _T_21 | _T_24; // @[LZD.scala 49:25]
  assign _T_26 = _T_13[0:0]; // @[LZD.scala 49:47]
  assign _T_27 = _T_20[0:0]; // @[LZD.scala 49:59]
  assign _T_28 = _T_21 ? _T_26 : _T_27; // @[LZD.scala 49:35]
  assign _T_30 = {_T_23,_T_25,_T_28}; // @[Cat.scala 29:58]
  assign _T_31 = ~ _T_30; // @[convert.scala 21:22]
  assign _T_32 = io_A[2:0]; // @[convert.scala 22:36]
  assign _T_33 = _T_31 < 3'h3; // @[Shift.scala 16:24]
  assign _T_34 = _T_31[1:0]; // @[Shift.scala 17:37]
  assign _T_35 = _T_34[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_32[0:0]; // @[Shift.scala 64:52]
  assign _T_38 = {_T_36,2'h0}; // @[Cat.scala 29:58]
  assign _T_39 = _T_35 ? _T_38 : _T_32; // @[Shift.scala 64:27]
  assign _T_40 = _T_34[0:0]; // @[Shift.scala 66:70]
  assign _T_42 = _T_39[1:0]; // @[Shift.scala 64:52]
  assign _T_43 = {_T_42,1'h0}; // @[Cat.scala 29:58]
  assign _T_44 = _T_40 ? _T_43 : _T_39; // @[Shift.scala 64:27]
  assign decA_fraction = _T_33 ? _T_44 : 3'h0; // @[Shift.scala 16:10]
  assign _T_48 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_50 = _T_3 ? _T_31 : _T_30; // @[convert.scala 25:42]
  assign _T_51 = {_T_48,_T_50}; // @[Cat.scala 29:58]
  assign _T_53 = io_A[4:0]; // @[convert.scala 29:56]
  assign _T_54 = _T_53 != 5'h0; // @[convert.scala 29:60]
  assign _T_55 = ~ _T_54; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_55; // @[convert.scala 29:39]
  assign _T_58 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_58 & _T_55; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_51); // @[convert.scala 32:24]
  assign _T_67 = io_B[5]; // @[convert.scala 18:24]
  assign _T_68 = io_B[4]; // @[convert.scala 18:40]
  assign _T_69 = _T_67 ^ _T_68; // @[convert.scala 18:36]
  assign _T_70 = io_B[4:1]; // @[convert.scala 19:24]
  assign _T_71 = io_B[3:0]; // @[convert.scala 19:43]
  assign _T_72 = _T_70 ^ _T_71; // @[convert.scala 19:39]
  assign _T_73 = _T_72[3:2]; // @[LZD.scala 43:32]
  assign _T_74 = _T_73 != 2'h0; // @[LZD.scala 39:14]
  assign _T_75 = _T_73[1]; // @[LZD.scala 39:21]
  assign _T_76 = _T_73[0]; // @[LZD.scala 39:30]
  assign _T_77 = ~ _T_76; // @[LZD.scala 39:27]
  assign _T_78 = _T_75 | _T_77; // @[LZD.scala 39:25]
  assign _T_79 = {_T_74,_T_78}; // @[Cat.scala 29:58]
  assign _T_80 = _T_72[1:0]; // @[LZD.scala 44:32]
  assign _T_81 = _T_80 != 2'h0; // @[LZD.scala 39:14]
  assign _T_82 = _T_80[1]; // @[LZD.scala 39:21]
  assign _T_83 = _T_80[0]; // @[LZD.scala 39:30]
  assign _T_84 = ~ _T_83; // @[LZD.scala 39:27]
  assign _T_85 = _T_82 | _T_84; // @[LZD.scala 39:25]
  assign _T_86 = {_T_81,_T_85}; // @[Cat.scala 29:58]
  assign _T_87 = _T_79[1]; // @[Shift.scala 12:21]
  assign _T_88 = _T_86[1]; // @[Shift.scala 12:21]
  assign _T_89 = _T_87 | _T_88; // @[LZD.scala 49:16]
  assign _T_90 = ~ _T_88; // @[LZD.scala 49:27]
  assign _T_91 = _T_87 | _T_90; // @[LZD.scala 49:25]
  assign _T_92 = _T_79[0:0]; // @[LZD.scala 49:47]
  assign _T_93 = _T_86[0:0]; // @[LZD.scala 49:59]
  assign _T_94 = _T_87 ? _T_92 : _T_93; // @[LZD.scala 49:35]
  assign _T_96 = {_T_89,_T_91,_T_94}; // @[Cat.scala 29:58]
  assign _T_97 = ~ _T_96; // @[convert.scala 21:22]
  assign _T_98 = io_B[2:0]; // @[convert.scala 22:36]
  assign _T_99 = _T_97 < 3'h3; // @[Shift.scala 16:24]
  assign _T_100 = _T_97[1:0]; // @[Shift.scala 17:37]
  assign _T_101 = _T_100[1]; // @[Shift.scala 12:21]
  assign _T_102 = _T_98[0:0]; // @[Shift.scala 64:52]
  assign _T_104 = {_T_102,2'h0}; // @[Cat.scala 29:58]
  assign _T_105 = _T_101 ? _T_104 : _T_98; // @[Shift.scala 64:27]
  assign _T_106 = _T_100[0:0]; // @[Shift.scala 66:70]
  assign _T_108 = _T_105[1:0]; // @[Shift.scala 64:52]
  assign _T_109 = {_T_108,1'h0}; // @[Cat.scala 29:58]
  assign _T_110 = _T_106 ? _T_109 : _T_105; // @[Shift.scala 64:27]
  assign decB_fraction = _T_99 ? _T_110 : 3'h0; // @[Shift.scala 16:10]
  assign _T_114 = _T_69 == 1'h0; // @[convert.scala 25:26]
  assign _T_116 = _T_69 ? _T_97 : _T_96; // @[convert.scala 25:42]
  assign _T_117 = {_T_114,_T_116}; // @[Cat.scala 29:58]
  assign _T_119 = io_B[4:0]; // @[convert.scala 29:56]
  assign _T_120 = _T_119 != 5'h0; // @[convert.scala 29:60]
  assign _T_121 = ~ _T_120; // @[convert.scala 29:41]
  assign decB_isNaR = _T_67 & _T_121; // @[convert.scala 29:39]
  assign _T_124 = _T_67 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_124 & _T_121; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_117); // @[convert.scala 32:24]
  assign _T_133 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_134 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_133,_T_134,decA_fraction,3'h0}; // @[Cat.scala 29:58]
  assign _T_137 = ~ _T_67; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_67,_T_137,decB_fraction,5'h0}; // @[Cat.scala 29:58]
  assign _T_140 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_140 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_141 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_142 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_143 = _T_142 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_144 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_145 = decA_isZero & _T_144; // @[PositDivisionSqrt.scala 94:43]
  assign _T_146 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_147 = _T_145 & _T_146; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_148 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_149 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_148 & _T_149; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_148 & _T_58; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_152 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_152; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 4'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_153 = sigX_Z[9]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_154 = sigX_Z[7]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_153 ^ _T_154; // @[PositDivisionSqrt.scala 113:50]
  assign _T_155 = cycleNum == 4'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_155 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_156 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_157 = _T_156 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_158 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_159 = entering & _T_158; // @[PositDivisionSqrt.scala 117:30]
  assign _T_161 = io_sqrtOp ? 4'h8 : 4'ha; // @[PositDivisionSqrt.scala 119:26]
  assign _T_162 = entering_normalCase ? _T_161 : 4'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{3'd0}, _T_159}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_163 = _GEN_9 | _T_162; // @[PositDivisionSqrt.scala 117:64]
  assign _T_165 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_166 = _T_156 & _T_165; // @[PositDivisionSqrt.scala 123:27]
  assign _T_168 = cycleNum - 4'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_169 = _T_166 ? _T_168 : 4'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _T_170 = _T_163 | _T_169; // @[PositDivisionSqrt.scala 122:64]
  assign _T_172 = _T_156 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_10 = {{3'd0}, _T_172}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_174 = _T_170 | _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  assign _T_175 = decA_scale[3:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_177 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_178 = entering_normalCase & _T_177; // @[PositDivisionSqrt.scala 137:28]
  assign _T_179 = 16'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign _T_180 = _T_179[15:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_181 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_182 = ready & _T_181; // @[PositDivisionSqrt.scala 148:23]
  assign _T_183 = _T_182 ? sigA_S : 10'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_184 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_185 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_186 = _T_185[9:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_187 = _T_184 ? _T_186 : 10'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_188 = _T_183 | _T_187; // @[PositDivisionSqrt.scala 148:66]
  assign _T_189 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_190 = _T_189 ? rem_Z : 10'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_188 | _T_190; // @[PositDivisionSqrt.scala 149:66]
  assign _T_192 = ready & _T_177; // @[PositDivisionSqrt.scala 152:29]
  assign _T_193 = _T_192 ? sigB_S : 10'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_194 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_195 = _T_194 ? 7'h40 : 7'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_11 = {{3'd0}, _T_195}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_196 = _T_193 | _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  assign _T_198 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_199 = _T_189 & _T_198; // @[PositDivisionSqrt.scala 154:30]
  assign _T_200 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_203 = {signB_Z,_T_200,fractB_Z,5'h0}; // @[Cat.scala 29:58]
  assign _T_204 = _T_199 ? _T_203 : 10'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_205 = _T_196 | _T_204; // @[PositDivisionSqrt.scala 153:93]
  assign _T_207 = _T_189 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_208 = rem[9:9]; // @[PositDivisionSqrt.scala 156:83]
  assign _T_210 = _T_208 ? 6'h3f : 6'h0; // @[Bitwise.scala 71:12]
  assign bitMask = _T_180[8:0]; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  assign _GEN_12 = {{3'd0}, _T_210}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_211 = bitMask & _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_13 = {{1'd0}, _T_211}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_212 = sigX_Z | _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  assign _T_213 = bitMask[8:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_14 = {{2'd0}, _T_213}; // @[PositDivisionSqrt.scala 156:89]
  assign _T_214 = _T_212 | _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  assign _T_215 = _T_207 ? _T_214 : 10'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_205 | _T_215; // @[PositDivisionSqrt.scala 154:93]
  assign _T_217 = trialTerm[9:9]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_218 = _T_208 ^ _T_217; // @[PositDivisionSqrt.scala 162:40]
  assign _T_221 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_223 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_224 = _T_218 ? _T_221 : _T_223; // @[PositDivisionSqrt.scala 161:92]
  assign _T_229 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_230 = _T_229[9:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_232 = _T_230 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_236 = _T_230 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_237 = _T_218 ? _T_232 : _T_236; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_224 : _T_237; // @[PositDivisionSqrt.scala 159:27]
  assign _T_238 = trialRem != 10'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_238 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_239 = rem != 10'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_239 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_241 = trialRem[9:9]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_242 = _T_217 ^ _T_241; // @[PositDivisionSqrt.scala 176:49]
  assign _T_243 = ~ _T_242; // @[PositDivisionSqrt.scala 176:29]
  assign _T_244 = sigX_Z[9:9]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_245 = ~ _T_244; // @[PositDivisionSqrt.scala 178:49]
  assign _T_247 = remIsZero ? _T_244 : _T_243; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_245 : _T_247; // @[Mux.scala 87:16]
  assign _T_248 = cycleNum > 4'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_249 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_250 = _T_248 & _T_249; // @[PositDivisionSqrt.scala 183:48]
  assign _T_251 = entering_normalCase | _T_250; // @[PositDivisionSqrt.scala 183:28]
  assign _T_254 = _T_189 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_255 = entering_normalCase | _T_254; // @[PositDivisionSqrt.scala 187:28]
  assign _T_258 = {newBit, 9'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_259 = _T_192 ? _T_258 : 10'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_261 = _T_194 ? 8'h80 : 8'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_15 = {{2'd0}, _T_261}; // @[PositDivisionSqrt.scala 188:78]
  assign _T_262 = _T_259 | _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  assign _GEN_16 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_264 = sigX_Z | _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  assign _T_265 = _T_189 ? _T_264 : 10'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_266 = _T_262 | _T_265; // @[PositDivisionSqrt.scala 189:78]
  assign _T_268 = {_T_244, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_268 : {{1'd0}, _T_244}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_17 = {{8'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  assign _T_271 = realSigX[6:4]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_272 = realSigX[5:3]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_271 : _T_272; // @[PositDivisionSqrt.scala 198:21]
  assign _T_273 = realSigX[9]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_274 = realSigX[7]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_275 = _T_273 ^ _T_274; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_275; // @[PositDivisionSqrt.scala 205:23]
  assign _T_277 = realSigX[6]; // @[PositDivisionSqrt.scala 206:56]
  assign notNeedSubTwo = _T_273 ^ _T_277; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_278 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_278; // @[PositDivisionSqrt.scala 208:36]
  assign _T_279 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_280 = {1'b0,$signed(_T_279)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_18 = {{2{_T_280[2]}},_T_280}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_282 = $signed(scale_Z) - $signed(_GEN_18); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_282); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-5'sh5); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(5'sh4); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[9:9]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_284 = underflow ? $signed(-5'sh5) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_285 = overflow ? $signed(5'sh4) : $signed(_T_284); // @[Mux.scala 87:16]
  assign _T_286 = realSigX[3:1]; // @[PositDivisionSqrt.scala 224:48]
  assign _T_287 = realSigX[2:0]; // @[PositDivisionSqrt.scala 224:64]
  assign decQ_grs = scaleNotChange ? _T_286 : _T_287; // @[PositDivisionSqrt.scala 224:23]
  assign outValid = cycleNum == 4'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_19 = _T_285[3:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_19); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_294 = decQ_scale[3:3]; // @[convert.scala 49:36]
  assign _T_296 = ~ decQ_scale; // @[convert.scala 50:36]
  assign _T_297 = $signed(_T_296); // @[convert.scala 50:36]
  assign _T_298 = _T_294 ? $signed(_T_297) : $signed(decQ_scale); // @[convert.scala 50:28]
  assign _T_299 = _T_294 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_300 = ~ _T_299; // @[convert.scala 53:34]
  assign _T_303 = {_T_300,_T_299,realFrac,decQ_grs}; // @[Cat.scala 29:58]
  assign _T_304 = $unsigned(_T_298); // @[Shift.scala 39:17]
  assign _T_305 = _T_304 < 4'h8; // @[Shift.scala 39:24]
  assign _T_306 = _T_298[2:0]; // @[Shift.scala 40:44]
  assign _T_307 = _T_303[7:4]; // @[Shift.scala 90:30]
  assign _T_308 = _T_303[3:0]; // @[Shift.scala 90:48]
  assign _T_309 = _T_308 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{3'd0}, _T_309}; // @[Shift.scala 90:39]
  assign _T_310 = _T_307 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_311 = _T_306[2]; // @[Shift.scala 12:21]
  assign _T_312 = _T_303[7]; // @[Shift.scala 12:21]
  assign _T_314 = _T_312 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_315 = {_T_314,_T_310}; // @[Cat.scala 29:58]
  assign _T_316 = _T_311 ? _T_315 : _T_303; // @[Shift.scala 91:22]
  assign _T_317 = _T_306[1:0]; // @[Shift.scala 92:77]
  assign _T_318 = _T_316[7:2]; // @[Shift.scala 90:30]
  assign _T_319 = _T_316[1:0]; // @[Shift.scala 90:48]
  assign _T_320 = _T_319 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{5'd0}, _T_320}; // @[Shift.scala 90:39]
  assign _T_321 = _T_318 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_322 = _T_317[1]; // @[Shift.scala 12:21]
  assign _T_323 = _T_316[7]; // @[Shift.scala 12:21]
  assign _T_325 = _T_323 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_326 = {_T_325,_T_321}; // @[Cat.scala 29:58]
  assign _T_327 = _T_322 ? _T_326 : _T_316; // @[Shift.scala 91:22]
  assign _T_328 = _T_317[0:0]; // @[Shift.scala 92:77]
  assign _T_329 = _T_327[7:1]; // @[Shift.scala 90:30]
  assign _T_330 = _T_327[0:0]; // @[Shift.scala 90:48]
  assign _GEN_22 = {{6'd0}, _T_330}; // @[Shift.scala 90:39]
  assign _T_332 = _T_329 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_334 = _T_327[7]; // @[Shift.scala 12:21]
  assign _T_335 = {_T_334,_T_332}; // @[Cat.scala 29:58]
  assign _T_336 = _T_328 ? _T_335 : _T_327; // @[Shift.scala 91:22]
  assign _T_339 = _T_312 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_340 = _T_305 ? _T_336 : _T_339; // @[Shift.scala 39:10]
  assign _T_341 = _T_340[3]; // @[convert.scala 55:31]
  assign _T_342 = _T_340[2]; // @[convert.scala 56:31]
  assign _T_343 = _T_340[1]; // @[convert.scala 57:31]
  assign _T_344 = _T_340[0]; // @[convert.scala 58:31]
  assign _T_345 = _T_340[7:3]; // @[convert.scala 59:69]
  assign _T_346 = _T_345 != 5'h0; // @[convert.scala 59:81]
  assign _T_347 = ~ _T_346; // @[convert.scala 59:50]
  assign _T_349 = _T_345 == 5'h1f; // @[convert.scala 60:81]
  assign _T_350 = _T_341 | _T_343; // @[convert.scala 61:44]
  assign _T_351 = _T_350 | _T_344; // @[convert.scala 61:52]
  assign _T_352 = _T_342 & _T_351; // @[convert.scala 61:36]
  assign _T_353 = ~ _T_349; // @[convert.scala 62:63]
  assign _T_354 = _T_353 & _T_352; // @[convert.scala 62:103]
  assign _T_355 = _T_347 | _T_354; // @[convert.scala 62:60]
  assign _GEN_23 = {{4'd0}, _T_355}; // @[convert.scala 63:56]
  assign _T_358 = _T_345 + _GEN_23; // @[convert.scala 63:56]
  assign _T_359 = {decQ_sign,_T_358}; // @[Cat.scala 29:58]
  assign _T_361 = isZero_Z ? 6'h0 : _T_359; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_198; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 6'h20 : _T_361; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 4'h0;
    end else begin
      if (_T_157) begin
        cycleNum <= _T_174;
      end
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_141;
      end else begin
        isNaR_Z <= _T_143;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_147;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_175[2]}},_T_175};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_178) begin
      signB_Z <= _T_67;
    end
    if (_T_178) begin
      if (_T_99) begin
        if (_T_106) begin
          fractB_Z <= _T_109;
        end else begin
          if (_T_101) begin
            fractB_Z <= _T_104;
          end else begin
            fractB_Z <= _T_98;
          end
        end
      end else begin
        fractB_Z <= 3'h0;
      end
    end
    if (_T_251) begin
      if (ready) begin
        if (_T_218) begin
          rem_Z <= _T_221;
        end else begin
          rem_Z <= _T_223;
        end
      end else begin
        if (_T_218) begin
          rem_Z <= _T_232;
        end else begin
          rem_Z <= _T_236;
        end
      end
    end
    if (_T_255) begin
      sigX_Z <= _T_266;
    end
  end
endmodule
