module PositMulDec4_0(
  input        clock,
  input        reset,
  input  [3:0] io_A,
  input  [3:0] io_B,
  output [2:0] io_sigA,
  output [2:0] io_sigB,
  output [2:0] io_decAscale,
  output [2:0] io_decBscale,
  output       io_decAisNar,
  output       io_decBisNar,
  output       io_decAisZero,
  output       io_decBisZero
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [1:0] _T_4; // @[convert.scala 19:24]
  wire [1:0] _T_5; // @[convert.scala 19:43]
  wire [1:0] _T_6; // @[convert.scala 19:39]
  wire  _T_7; // @[LZD.scala 39:14]
  wire  _T_8; // @[LZD.scala 39:21]
  wire  _T_9; // @[LZD.scala 39:30]
  wire  _T_10; // @[LZD.scala 39:27]
  wire  _T_11; // @[LZD.scala 39:25]
  wire [1:0] _T_12; // @[Cat.scala 29:58]
  wire [1:0] _T_13; // @[convert.scala 21:22]
  wire  _T_14; // @[convert.scala 22:36]
  wire  _T_15; // @[Shift.scala 16:24]
  wire  _T_16; // @[Shift.scala 17:37]
  wire  _T_18; // @[Shift.scala 63:39]
  wire  decA_fraction; // @[Shift.scala 16:10]
  wire  _T_22; // @[convert.scala 25:26]
  wire [1:0] _T_24; // @[convert.scala 25:42]
  wire [2:0] _T_25; // @[Cat.scala 29:58]
  wire [2:0] _T_27; // @[convert.scala 29:56]
  wire  _T_28; // @[convert.scala 29:60]
  wire  _T_29; // @[convert.scala 29:41]
  wire  _T_32; // @[convert.scala 30:19]
  wire  _T_41; // @[convert.scala 18:24]
  wire  _T_42; // @[convert.scala 18:40]
  wire  _T_43; // @[convert.scala 18:36]
  wire [1:0] _T_44; // @[convert.scala 19:24]
  wire [1:0] _T_45; // @[convert.scala 19:43]
  wire [1:0] _T_46; // @[convert.scala 19:39]
  wire  _T_47; // @[LZD.scala 39:14]
  wire  _T_48; // @[LZD.scala 39:21]
  wire  _T_49; // @[LZD.scala 39:30]
  wire  _T_50; // @[LZD.scala 39:27]
  wire  _T_51; // @[LZD.scala 39:25]
  wire [1:0] _T_52; // @[Cat.scala 29:58]
  wire [1:0] _T_53; // @[convert.scala 21:22]
  wire  _T_54; // @[convert.scala 22:36]
  wire  _T_55; // @[Shift.scala 16:24]
  wire  _T_56; // @[Shift.scala 17:37]
  wire  _T_58; // @[Shift.scala 63:39]
  wire  decB_fraction; // @[Shift.scala 16:10]
  wire  _T_62; // @[convert.scala 25:26]
  wire [1:0] _T_64; // @[convert.scala 25:42]
  wire [2:0] _T_65; // @[Cat.scala 29:58]
  wire [2:0] _T_67; // @[convert.scala 29:56]
  wire  _T_68; // @[convert.scala 29:60]
  wire  _T_69; // @[convert.scala 29:41]
  wire  _T_72; // @[convert.scala 30:19]
  wire  _T_80; // @[PositMulDec.scala 31:34]
  wire [2:0] _T_82; // @[Cat.scala 29:58]
  wire  _T_84; // @[PositMulDec.scala 32:34]
  wire [2:0] _T_86; // @[Cat.scala 29:58]
  assign _T_1 = io_A[3]; // @[convert.scala 18:24]
  assign _T_2 = io_A[2]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[2:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[1:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6 != 2'h0; // @[LZD.scala 39:14]
  assign _T_8 = _T_6[1]; // @[LZD.scala 39:21]
  assign _T_9 = _T_6[0]; // @[LZD.scala 39:30]
  assign _T_10 = ~ _T_9; // @[LZD.scala 39:27]
  assign _T_11 = _T_8 | _T_10; // @[LZD.scala 39:25]
  assign _T_12 = {_T_7,_T_11}; // @[Cat.scala 29:58]
  assign _T_13 = ~ _T_12; // @[convert.scala 21:22]
  assign _T_14 = io_A[0:0]; // @[convert.scala 22:36]
  assign _T_15 = _T_13 < 2'h1; // @[Shift.scala 16:24]
  assign _T_16 = _T_13[0]; // @[Shift.scala 17:37]
  assign _T_18 = _T_16 ? 1'h0 : _T_14; // @[Shift.scala 63:39]
  assign decA_fraction = _T_15 & _T_18; // @[Shift.scala 16:10]
  assign _T_22 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_24 = _T_3 ? _T_13 : _T_12; // @[convert.scala 25:42]
  assign _T_25 = {_T_22,_T_24}; // @[Cat.scala 29:58]
  assign _T_27 = io_A[2:0]; // @[convert.scala 29:56]
  assign _T_28 = _T_27 != 3'h0; // @[convert.scala 29:60]
  assign _T_29 = ~ _T_28; // @[convert.scala 29:41]
  assign _T_32 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign _T_41 = io_B[3]; // @[convert.scala 18:24]
  assign _T_42 = io_B[2]; // @[convert.scala 18:40]
  assign _T_43 = _T_41 ^ _T_42; // @[convert.scala 18:36]
  assign _T_44 = io_B[2:1]; // @[convert.scala 19:24]
  assign _T_45 = io_B[1:0]; // @[convert.scala 19:43]
  assign _T_46 = _T_44 ^ _T_45; // @[convert.scala 19:39]
  assign _T_47 = _T_46 != 2'h0; // @[LZD.scala 39:14]
  assign _T_48 = _T_46[1]; // @[LZD.scala 39:21]
  assign _T_49 = _T_46[0]; // @[LZD.scala 39:30]
  assign _T_50 = ~ _T_49; // @[LZD.scala 39:27]
  assign _T_51 = _T_48 | _T_50; // @[LZD.scala 39:25]
  assign _T_52 = {_T_47,_T_51}; // @[Cat.scala 29:58]
  assign _T_53 = ~ _T_52; // @[convert.scala 21:22]
  assign _T_54 = io_B[0:0]; // @[convert.scala 22:36]
  assign _T_55 = _T_53 < 2'h1; // @[Shift.scala 16:24]
  assign _T_56 = _T_53[0]; // @[Shift.scala 17:37]
  assign _T_58 = _T_56 ? 1'h0 : _T_54; // @[Shift.scala 63:39]
  assign decB_fraction = _T_55 & _T_58; // @[Shift.scala 16:10]
  assign _T_62 = _T_43 == 1'h0; // @[convert.scala 25:26]
  assign _T_64 = _T_43 ? _T_53 : _T_52; // @[convert.scala 25:42]
  assign _T_65 = {_T_62,_T_64}; // @[Cat.scala 29:58]
  assign _T_67 = io_B[2:0]; // @[convert.scala 29:56]
  assign _T_68 = _T_67 != 3'h0; // @[convert.scala 29:60]
  assign _T_69 = ~ _T_68; // @[convert.scala 29:41]
  assign _T_72 = _T_41 == 1'h0; // @[convert.scala 30:19]
  assign _T_80 = ~ _T_1; // @[PositMulDec.scala 31:34]
  assign _T_82 = {_T_1,_T_80,decA_fraction}; // @[Cat.scala 29:58]
  assign _T_84 = ~ _T_41; // @[PositMulDec.scala 32:34]
  assign _T_86 = {_T_41,_T_84,decB_fraction}; // @[Cat.scala 29:58]
  assign io_sigA = $signed(_T_82); // @[PositMulDec.scala 31:16]
  assign io_sigB = $signed(_T_86); // @[PositMulDec.scala 32:16]
  assign io_decAscale = $signed(_T_25); // @[PositMulDec.scala 33:16]
  assign io_decBscale = $signed(_T_65); // @[PositMulDec.scala 34:16]
  assign io_decAisNar = _T_1 & _T_29; // @[PositMulDec.scala 35:16]
  assign io_decBisNar = _T_41 & _T_69; // @[PositMulDec.scala 36:16]
  assign io_decAisZero = _T_32 & _T_29; // @[PositMulDec.scala 37:17]
  assign io_decBisZero = _T_72 & _T_69; // @[PositMulDec.scala 38:17]
endmodule
