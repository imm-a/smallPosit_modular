module FMA_Dec5_0(
  input        clock,
  input        reset,
  input  [4:0] io_A,
  input  [4:0] io_B,
  input  [4:0] io_C,
  output [3:0] io_sigA,
  output [3:0] io_sigB,
  output       io_outIsNaR,
  output       io_Csign,
  output       io_CisNar,
  output       io_CisZero,
  output [1:0] io_Cfrac,
  output [2:0] io_Ascale,
  output [2:0] io_Bscale,
  output [2:0] io_Cscale
);
  wire [5:0] _T_2; // @[FMA_Dec.scala 38:46]
  wire [4:0] realA; // @[FMA_Dec.scala 38:46]
  wire [5:0] _T_5; // @[FMA_Dec.scala 39:46]
  wire [4:0] realC; // @[FMA_Dec.scala 39:46]
  wire  _T_7; // @[convert.scala 18:24]
  wire  _T_8; // @[convert.scala 18:40]
  wire  _T_9; // @[convert.scala 18:36]
  wire [2:0] _T_10; // @[convert.scala 19:24]
  wire [2:0] _T_11; // @[convert.scala 19:43]
  wire [2:0] _T_12; // @[convert.scala 19:39]
  wire [1:0] _T_13; // @[LZD.scala 43:32]
  wire  _T_14; // @[LZD.scala 39:14]
  wire  _T_15; // @[LZD.scala 39:21]
  wire  _T_16; // @[LZD.scala 39:30]
  wire  _T_17; // @[LZD.scala 39:27]
  wire  _T_18; // @[LZD.scala 39:25]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  _T_20; // @[LZD.scala 44:32]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_24; // @[LZD.scala 55:32]
  wire  _T_25; // @[LZD.scala 55:20]
  wire [1:0] _T_26; // @[Cat.scala 29:58]
  wire [1:0] _T_27; // @[convert.scala 21:22]
  wire [1:0] _T_28; // @[convert.scala 22:36]
  wire  _T_29; // @[Shift.scala 16:24]
  wire  _T_30; // @[Shift.scala 17:37]
  wire  _T_32; // @[Shift.scala 64:52]
  wire [1:0] _T_33; // @[Cat.scala 29:58]
  wire [1:0] _T_34; // @[Shift.scala 64:27]
  wire [1:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_38; // @[convert.scala 25:26]
  wire [1:0] _T_40; // @[convert.scala 25:42]
  wire [2:0] _T_41; // @[Cat.scala 29:58]
  wire [3:0] _T_43; // @[convert.scala 29:56]
  wire  _T_44; // @[convert.scala 29:60]
  wire  _T_45; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_48; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire  _T_57; // @[convert.scala 18:24]
  wire  _T_58; // @[convert.scala 18:40]
  wire  _T_59; // @[convert.scala 18:36]
  wire [2:0] _T_60; // @[convert.scala 19:24]
  wire [2:0] _T_61; // @[convert.scala 19:43]
  wire [2:0] _T_62; // @[convert.scala 19:39]
  wire [1:0] _T_63; // @[LZD.scala 43:32]
  wire  _T_64; // @[LZD.scala 39:14]
  wire  _T_65; // @[LZD.scala 39:21]
  wire  _T_66; // @[LZD.scala 39:30]
  wire  _T_67; // @[LZD.scala 39:27]
  wire  _T_68; // @[LZD.scala 39:25]
  wire [1:0] _T_69; // @[Cat.scala 29:58]
  wire  _T_70; // @[LZD.scala 44:32]
  wire  _T_72; // @[Shift.scala 12:21]
  wire  _T_74; // @[LZD.scala 55:32]
  wire  _T_75; // @[LZD.scala 55:20]
  wire [1:0] _T_76; // @[Cat.scala 29:58]
  wire [1:0] _T_77; // @[convert.scala 21:22]
  wire [1:0] _T_78; // @[convert.scala 22:36]
  wire  _T_79; // @[Shift.scala 16:24]
  wire  _T_80; // @[Shift.scala 17:37]
  wire  _T_82; // @[Shift.scala 64:52]
  wire [1:0] _T_83; // @[Cat.scala 29:58]
  wire [1:0] _T_84; // @[Shift.scala 64:27]
  wire [1:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_88; // @[convert.scala 25:26]
  wire [1:0] _T_90; // @[convert.scala 25:42]
  wire [2:0] _T_91; // @[Cat.scala 29:58]
  wire [3:0] _T_93; // @[convert.scala 29:56]
  wire  _T_94; // @[convert.scala 29:60]
  wire  _T_95; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_98; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire  _T_107; // @[convert.scala 18:24]
  wire  _T_108; // @[convert.scala 18:40]
  wire  _T_109; // @[convert.scala 18:36]
  wire [2:0] _T_110; // @[convert.scala 19:24]
  wire [2:0] _T_111; // @[convert.scala 19:43]
  wire [2:0] _T_112; // @[convert.scala 19:39]
  wire [1:0] _T_113; // @[LZD.scala 43:32]
  wire  _T_114; // @[LZD.scala 39:14]
  wire  _T_115; // @[LZD.scala 39:21]
  wire  _T_116; // @[LZD.scala 39:30]
  wire  _T_117; // @[LZD.scala 39:27]
  wire  _T_118; // @[LZD.scala 39:25]
  wire [1:0] _T_119; // @[Cat.scala 29:58]
  wire  _T_120; // @[LZD.scala 44:32]
  wire  _T_122; // @[Shift.scala 12:21]
  wire  _T_124; // @[LZD.scala 55:32]
  wire  _T_125; // @[LZD.scala 55:20]
  wire [1:0] _T_126; // @[Cat.scala 29:58]
  wire [1:0] _T_127; // @[convert.scala 21:22]
  wire [1:0] _T_128; // @[convert.scala 22:36]
  wire  _T_129; // @[Shift.scala 16:24]
  wire  _T_130; // @[Shift.scala 17:37]
  wire  _T_132; // @[Shift.scala 64:52]
  wire [1:0] _T_133; // @[Cat.scala 29:58]
  wire [1:0] _T_134; // @[Shift.scala 64:27]
  wire  _T_138; // @[convert.scala 25:26]
  wire [1:0] _T_140; // @[convert.scala 25:42]
  wire [2:0] _T_141; // @[Cat.scala 29:58]
  wire [3:0] _T_143; // @[convert.scala 29:56]
  wire  _T_144; // @[convert.scala 29:60]
  wire  _T_145; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_148; // @[convert.scala 30:19]
  wire  _T_156; // @[FMA_Dec.scala 46:30]
  wire  _T_158; // @[FMA_Dec.scala 49:34]
  wire  _T_159; // @[FMA_Dec.scala 49:47]
  wire  _T_160; // @[FMA_Dec.scala 49:45]
  wire [3:0] _T_162; // @[Cat.scala 29:58]
  wire  _T_164; // @[FMA_Dec.scala 50:34]
  wire  _T_165; // @[FMA_Dec.scala 50:47]
  wire  _T_166; // @[FMA_Dec.scala 50:45]
  wire [3:0] _T_168; // @[Cat.scala 29:58]
  assign _T_2 = {{1'd0}, io_A}; // @[FMA_Dec.scala 38:46]
  assign realA = _T_2[4:0]; // @[FMA_Dec.scala 38:46]
  assign _T_5 = {{1'd0}, io_C}; // @[FMA_Dec.scala 39:46]
  assign realC = _T_5[4:0]; // @[FMA_Dec.scala 39:46]
  assign _T_7 = realA[4]; // @[convert.scala 18:24]
  assign _T_8 = realA[3]; // @[convert.scala 18:40]
  assign _T_9 = _T_7 ^ _T_8; // @[convert.scala 18:36]
  assign _T_10 = realA[3:1]; // @[convert.scala 19:24]
  assign _T_11 = realA[2:0]; // @[convert.scala 19:43]
  assign _T_12 = _T_10 ^ _T_11; // @[convert.scala 19:39]
  assign _T_13 = _T_12[2:1]; // @[LZD.scala 43:32]
  assign _T_14 = _T_13 != 2'h0; // @[LZD.scala 39:14]
  assign _T_15 = _T_13[1]; // @[LZD.scala 39:21]
  assign _T_16 = _T_13[0]; // @[LZD.scala 39:30]
  assign _T_17 = ~ _T_16; // @[LZD.scala 39:27]
  assign _T_18 = _T_15 | _T_17; // @[LZD.scala 39:25]
  assign _T_19 = {_T_14,_T_18}; // @[Cat.scala 29:58]
  assign _T_20 = _T_12[0:0]; // @[LZD.scala 44:32]
  assign _T_22 = _T_19[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_19[0:0]; // @[LZD.scala 55:32]
  assign _T_25 = _T_22 ? _T_24 : _T_20; // @[LZD.scala 55:20]
  assign _T_26 = {_T_22,_T_25}; // @[Cat.scala 29:58]
  assign _T_27 = ~ _T_26; // @[convert.scala 21:22]
  assign _T_28 = realA[1:0]; // @[convert.scala 22:36]
  assign _T_29 = _T_27 < 2'h2; // @[Shift.scala 16:24]
  assign _T_30 = _T_27[0]; // @[Shift.scala 17:37]
  assign _T_32 = _T_28[0:0]; // @[Shift.scala 64:52]
  assign _T_33 = {_T_32,1'h0}; // @[Cat.scala 29:58]
  assign _T_34 = _T_30 ? _T_33 : _T_28; // @[Shift.scala 64:27]
  assign decA_fraction = _T_29 ? _T_34 : 2'h0; // @[Shift.scala 16:10]
  assign _T_38 = _T_9 == 1'h0; // @[convert.scala 25:26]
  assign _T_40 = _T_9 ? _T_27 : _T_26; // @[convert.scala 25:42]
  assign _T_41 = {_T_38,_T_40}; // @[Cat.scala 29:58]
  assign _T_43 = realA[3:0]; // @[convert.scala 29:56]
  assign _T_44 = _T_43 != 4'h0; // @[convert.scala 29:60]
  assign _T_45 = ~ _T_44; // @[convert.scala 29:41]
  assign decA_isNaR = _T_7 & _T_45; // @[convert.scala 29:39]
  assign _T_48 = _T_7 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_48 & _T_45; // @[convert.scala 30:41]
  assign _T_57 = io_B[4]; // @[convert.scala 18:24]
  assign _T_58 = io_B[3]; // @[convert.scala 18:40]
  assign _T_59 = _T_57 ^ _T_58; // @[convert.scala 18:36]
  assign _T_60 = io_B[3:1]; // @[convert.scala 19:24]
  assign _T_61 = io_B[2:0]; // @[convert.scala 19:43]
  assign _T_62 = _T_60 ^ _T_61; // @[convert.scala 19:39]
  assign _T_63 = _T_62[2:1]; // @[LZD.scala 43:32]
  assign _T_64 = _T_63 != 2'h0; // @[LZD.scala 39:14]
  assign _T_65 = _T_63[1]; // @[LZD.scala 39:21]
  assign _T_66 = _T_63[0]; // @[LZD.scala 39:30]
  assign _T_67 = ~ _T_66; // @[LZD.scala 39:27]
  assign _T_68 = _T_65 | _T_67; // @[LZD.scala 39:25]
  assign _T_69 = {_T_64,_T_68}; // @[Cat.scala 29:58]
  assign _T_70 = _T_62[0:0]; // @[LZD.scala 44:32]
  assign _T_72 = _T_69[1]; // @[Shift.scala 12:21]
  assign _T_74 = _T_69[0:0]; // @[LZD.scala 55:32]
  assign _T_75 = _T_72 ? _T_74 : _T_70; // @[LZD.scala 55:20]
  assign _T_76 = {_T_72,_T_75}; // @[Cat.scala 29:58]
  assign _T_77 = ~ _T_76; // @[convert.scala 21:22]
  assign _T_78 = io_B[1:0]; // @[convert.scala 22:36]
  assign _T_79 = _T_77 < 2'h2; // @[Shift.scala 16:24]
  assign _T_80 = _T_77[0]; // @[Shift.scala 17:37]
  assign _T_82 = _T_78[0:0]; // @[Shift.scala 64:52]
  assign _T_83 = {_T_82,1'h0}; // @[Cat.scala 29:58]
  assign _T_84 = _T_80 ? _T_83 : _T_78; // @[Shift.scala 64:27]
  assign decB_fraction = _T_79 ? _T_84 : 2'h0; // @[Shift.scala 16:10]
  assign _T_88 = _T_59 == 1'h0; // @[convert.scala 25:26]
  assign _T_90 = _T_59 ? _T_77 : _T_76; // @[convert.scala 25:42]
  assign _T_91 = {_T_88,_T_90}; // @[Cat.scala 29:58]
  assign _T_93 = io_B[3:0]; // @[convert.scala 29:56]
  assign _T_94 = _T_93 != 4'h0; // @[convert.scala 29:60]
  assign _T_95 = ~ _T_94; // @[convert.scala 29:41]
  assign decB_isNaR = _T_57 & _T_95; // @[convert.scala 29:39]
  assign _T_98 = _T_57 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_98 & _T_95; // @[convert.scala 30:41]
  assign _T_107 = realC[4]; // @[convert.scala 18:24]
  assign _T_108 = realC[3]; // @[convert.scala 18:40]
  assign _T_109 = _T_107 ^ _T_108; // @[convert.scala 18:36]
  assign _T_110 = realC[3:1]; // @[convert.scala 19:24]
  assign _T_111 = realC[2:0]; // @[convert.scala 19:43]
  assign _T_112 = _T_110 ^ _T_111; // @[convert.scala 19:39]
  assign _T_113 = _T_112[2:1]; // @[LZD.scala 43:32]
  assign _T_114 = _T_113 != 2'h0; // @[LZD.scala 39:14]
  assign _T_115 = _T_113[1]; // @[LZD.scala 39:21]
  assign _T_116 = _T_113[0]; // @[LZD.scala 39:30]
  assign _T_117 = ~ _T_116; // @[LZD.scala 39:27]
  assign _T_118 = _T_115 | _T_117; // @[LZD.scala 39:25]
  assign _T_119 = {_T_114,_T_118}; // @[Cat.scala 29:58]
  assign _T_120 = _T_112[0:0]; // @[LZD.scala 44:32]
  assign _T_122 = _T_119[1]; // @[Shift.scala 12:21]
  assign _T_124 = _T_119[0:0]; // @[LZD.scala 55:32]
  assign _T_125 = _T_122 ? _T_124 : _T_120; // @[LZD.scala 55:20]
  assign _T_126 = {_T_122,_T_125}; // @[Cat.scala 29:58]
  assign _T_127 = ~ _T_126; // @[convert.scala 21:22]
  assign _T_128 = realC[1:0]; // @[convert.scala 22:36]
  assign _T_129 = _T_127 < 2'h2; // @[Shift.scala 16:24]
  assign _T_130 = _T_127[0]; // @[Shift.scala 17:37]
  assign _T_132 = _T_128[0:0]; // @[Shift.scala 64:52]
  assign _T_133 = {_T_132,1'h0}; // @[Cat.scala 29:58]
  assign _T_134 = _T_130 ? _T_133 : _T_128; // @[Shift.scala 64:27]
  assign _T_138 = _T_109 == 1'h0; // @[convert.scala 25:26]
  assign _T_140 = _T_109 ? _T_127 : _T_126; // @[convert.scala 25:42]
  assign _T_141 = {_T_138,_T_140}; // @[Cat.scala 29:58]
  assign _T_143 = realC[3:0]; // @[convert.scala 29:56]
  assign _T_144 = _T_143 != 4'h0; // @[convert.scala 29:60]
  assign _T_145 = ~ _T_144; // @[convert.scala 29:41]
  assign decC_isNaR = _T_107 & _T_145; // @[convert.scala 29:39]
  assign _T_148 = _T_107 == 1'h0; // @[convert.scala 30:19]
  assign _T_156 = decA_isNaR | decB_isNaR; // @[FMA_Dec.scala 46:30]
  assign _T_158 = ~ _T_7; // @[FMA_Dec.scala 49:34]
  assign _T_159 = ~ decA_isZero; // @[FMA_Dec.scala 49:47]
  assign _T_160 = _T_158 & _T_159; // @[FMA_Dec.scala 49:45]
  assign _T_162 = {_T_7,_T_160,decA_fraction}; // @[Cat.scala 29:58]
  assign _T_164 = ~ _T_57; // @[FMA_Dec.scala 50:34]
  assign _T_165 = ~ decB_isZero; // @[FMA_Dec.scala 50:47]
  assign _T_166 = _T_164 & _T_165; // @[FMA_Dec.scala 50:45]
  assign _T_168 = {_T_57,_T_166,decB_fraction}; // @[Cat.scala 29:58]
  assign io_sigA = $signed(_T_162); // @[FMA_Dec.scala 49:16]
  assign io_sigB = $signed(_T_168); // @[FMA_Dec.scala 50:16]
  assign io_outIsNaR = _T_156 | decC_isNaR; // @[FMA_Dec.scala 46:16]
  assign io_Csign = realC[4]; // @[FMA_Dec.scala 55:12]
  assign io_CisNar = _T_107 & _T_145; // @[FMA_Dec.scala 51:17]
  assign io_CisZero = _T_148 & _T_145; // @[FMA_Dec.scala 52:17]
  assign io_Cfrac = _T_129 ? _T_134 : 2'h0; // @[FMA_Dec.scala 53:17]
  assign io_Ascale = $signed(_T_41); // @[FMA_Dec.scala 47:13]
  assign io_Bscale = $signed(_T_91); // @[FMA_Dec.scala 48:13]
  assign io_Cscale = $signed(_T_141); // @[FMA_Dec.scala 54:16]
endmodule
