module PositFMA6_2(
  input        clock,
  input        reset,
  input        io_inValid,
  input  [1:0] io_fmaOp,
  input  [5:0] io_A,
  input  [5:0] io_B,
  input  [5:0] io_C,
  output [5:0] io_F,
  output       io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [5:0] _T_2; // @[Bitwise.scala 71:12]
  wire [5:0] _T_3; // @[PositFMA.scala 47:41]
  wire [5:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [5:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [5:0] _T_8; // @[Bitwise.scala 71:12]
  wire [5:0] _T_9; // @[PositFMA.scala 48:41]
  wire [5:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [5:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [3:0] _T_16; // @[convert.scala 19:24]
  wire [3:0] _T_17; // @[convert.scala 19:43]
  wire [3:0] _T_18; // @[convert.scala 19:39]
  wire [1:0] _T_19; // @[LZD.scala 43:32]
  wire  _T_20; // @[LZD.scala 39:14]
  wire  _T_21; // @[LZD.scala 39:21]
  wire  _T_22; // @[LZD.scala 39:30]
  wire  _T_23; // @[LZD.scala 39:27]
  wire  _T_24; // @[LZD.scala 39:25]
  wire [1:0] _T_25; // @[Cat.scala 29:58]
  wire [1:0] _T_26; // @[LZD.scala 44:32]
  wire  _T_27; // @[LZD.scala 39:14]
  wire  _T_28; // @[LZD.scala 39:21]
  wire  _T_29; // @[LZD.scala 39:30]
  wire  _T_30; // @[LZD.scala 39:27]
  wire  _T_31; // @[LZD.scala 39:25]
  wire [1:0] _T_32; // @[Cat.scala 29:58]
  wire  _T_33; // @[Shift.scala 12:21]
  wire  _T_34; // @[Shift.scala 12:21]
  wire  _T_35; // @[LZD.scala 49:16]
  wire  _T_36; // @[LZD.scala 49:27]
  wire  _T_37; // @[LZD.scala 49:25]
  wire  _T_38; // @[LZD.scala 49:47]
  wire  _T_39; // @[LZD.scala 49:59]
  wire  _T_40; // @[LZD.scala 49:35]
  wire [2:0] _T_42; // @[Cat.scala 29:58]
  wire [2:0] _T_43; // @[convert.scala 21:22]
  wire [2:0] _T_44; // @[convert.scala 22:36]
  wire  _T_45; // @[Shift.scala 16:24]
  wire [1:0] _T_46; // @[Shift.scala 17:37]
  wire  _T_47; // @[Shift.scala 12:21]
  wire  _T_48; // @[Shift.scala 64:52]
  wire [2:0] _T_50; // @[Cat.scala 29:58]
  wire [2:0] _T_51; // @[Shift.scala 64:27]
  wire  _T_52; // @[Shift.scala 66:70]
  wire [1:0] _T_54; // @[Shift.scala 64:52]
  wire [2:0] _T_55; // @[Cat.scala 29:58]
  wire [2:0] _T_56; // @[Shift.scala 64:27]
  wire [2:0] _T_57; // @[Shift.scala 16:10]
  wire [1:0] _T_58; // @[convert.scala 23:34]
  wire  decA_fraction; // @[convert.scala 24:34]
  wire  _T_60; // @[convert.scala 25:26]
  wire [2:0] _T_62; // @[convert.scala 25:42]
  wire [1:0] _T_65; // @[convert.scala 26:67]
  wire [1:0] _T_66; // @[convert.scala 26:51]
  wire [5:0] _T_67; // @[Cat.scala 29:58]
  wire [4:0] _T_69; // @[convert.scala 29:56]
  wire  _T_70; // @[convert.scala 29:60]
  wire  _T_71; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_74; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_83; // @[convert.scala 18:24]
  wire  _T_84; // @[convert.scala 18:40]
  wire  _T_85; // @[convert.scala 18:36]
  wire [3:0] _T_86; // @[convert.scala 19:24]
  wire [3:0] _T_87; // @[convert.scala 19:43]
  wire [3:0] _T_88; // @[convert.scala 19:39]
  wire [1:0] _T_89; // @[LZD.scala 43:32]
  wire  _T_90; // @[LZD.scala 39:14]
  wire  _T_91; // @[LZD.scala 39:21]
  wire  _T_92; // @[LZD.scala 39:30]
  wire  _T_93; // @[LZD.scala 39:27]
  wire  _T_94; // @[LZD.scala 39:25]
  wire [1:0] _T_95; // @[Cat.scala 29:58]
  wire [1:0] _T_96; // @[LZD.scala 44:32]
  wire  _T_97; // @[LZD.scala 39:14]
  wire  _T_98; // @[LZD.scala 39:21]
  wire  _T_99; // @[LZD.scala 39:30]
  wire  _T_100; // @[LZD.scala 39:27]
  wire  _T_101; // @[LZD.scala 39:25]
  wire [1:0] _T_102; // @[Cat.scala 29:58]
  wire  _T_103; // @[Shift.scala 12:21]
  wire  _T_104; // @[Shift.scala 12:21]
  wire  _T_105; // @[LZD.scala 49:16]
  wire  _T_106; // @[LZD.scala 49:27]
  wire  _T_107; // @[LZD.scala 49:25]
  wire  _T_108; // @[LZD.scala 49:47]
  wire  _T_109; // @[LZD.scala 49:59]
  wire  _T_110; // @[LZD.scala 49:35]
  wire [2:0] _T_112; // @[Cat.scala 29:58]
  wire [2:0] _T_113; // @[convert.scala 21:22]
  wire [2:0] _T_114; // @[convert.scala 22:36]
  wire  _T_115; // @[Shift.scala 16:24]
  wire [1:0] _T_116; // @[Shift.scala 17:37]
  wire  _T_117; // @[Shift.scala 12:21]
  wire  _T_118; // @[Shift.scala 64:52]
  wire [2:0] _T_120; // @[Cat.scala 29:58]
  wire [2:0] _T_121; // @[Shift.scala 64:27]
  wire  _T_122; // @[Shift.scala 66:70]
  wire [1:0] _T_124; // @[Shift.scala 64:52]
  wire [2:0] _T_125; // @[Cat.scala 29:58]
  wire [2:0] _T_126; // @[Shift.scala 64:27]
  wire [2:0] _T_127; // @[Shift.scala 16:10]
  wire [1:0] _T_128; // @[convert.scala 23:34]
  wire  decB_fraction; // @[convert.scala 24:34]
  wire  _T_130; // @[convert.scala 25:26]
  wire [2:0] _T_132; // @[convert.scala 25:42]
  wire [1:0] _T_135; // @[convert.scala 26:67]
  wire [1:0] _T_136; // @[convert.scala 26:51]
  wire [5:0] _T_137; // @[Cat.scala 29:58]
  wire [4:0] _T_139; // @[convert.scala 29:56]
  wire  _T_140; // @[convert.scala 29:60]
  wire  _T_141; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_144; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_153; // @[convert.scala 18:24]
  wire  _T_154; // @[convert.scala 18:40]
  wire  _T_155; // @[convert.scala 18:36]
  wire [3:0] _T_156; // @[convert.scala 19:24]
  wire [3:0] _T_157; // @[convert.scala 19:43]
  wire [3:0] _T_158; // @[convert.scala 19:39]
  wire [1:0] _T_159; // @[LZD.scala 43:32]
  wire  _T_160; // @[LZD.scala 39:14]
  wire  _T_161; // @[LZD.scala 39:21]
  wire  _T_162; // @[LZD.scala 39:30]
  wire  _T_163; // @[LZD.scala 39:27]
  wire  _T_164; // @[LZD.scala 39:25]
  wire [1:0] _T_165; // @[Cat.scala 29:58]
  wire [1:0] _T_166; // @[LZD.scala 44:32]
  wire  _T_167; // @[LZD.scala 39:14]
  wire  _T_168; // @[LZD.scala 39:21]
  wire  _T_169; // @[LZD.scala 39:30]
  wire  _T_170; // @[LZD.scala 39:27]
  wire  _T_171; // @[LZD.scala 39:25]
  wire [1:0] _T_172; // @[Cat.scala 29:58]
  wire  _T_173; // @[Shift.scala 12:21]
  wire  _T_174; // @[Shift.scala 12:21]
  wire  _T_175; // @[LZD.scala 49:16]
  wire  _T_176; // @[LZD.scala 49:27]
  wire  _T_177; // @[LZD.scala 49:25]
  wire  _T_178; // @[LZD.scala 49:47]
  wire  _T_179; // @[LZD.scala 49:59]
  wire  _T_180; // @[LZD.scala 49:35]
  wire [2:0] _T_182; // @[Cat.scala 29:58]
  wire [2:0] _T_183; // @[convert.scala 21:22]
  wire [2:0] _T_184; // @[convert.scala 22:36]
  wire  _T_185; // @[Shift.scala 16:24]
  wire [1:0] _T_186; // @[Shift.scala 17:37]
  wire  _T_187; // @[Shift.scala 12:21]
  wire  _T_188; // @[Shift.scala 64:52]
  wire [2:0] _T_190; // @[Cat.scala 29:58]
  wire [2:0] _T_191; // @[Shift.scala 64:27]
  wire  _T_192; // @[Shift.scala 66:70]
  wire [1:0] _T_194; // @[Shift.scala 64:52]
  wire [2:0] _T_195; // @[Cat.scala 29:58]
  wire [2:0] _T_196; // @[Shift.scala 64:27]
  wire [2:0] _T_197; // @[Shift.scala 16:10]
  wire [1:0] _T_198; // @[convert.scala 23:34]
  wire  decC_fraction; // @[convert.scala 24:34]
  wire  _T_200; // @[convert.scala 25:26]
  wire [2:0] _T_202; // @[convert.scala 25:42]
  wire [1:0] _T_205; // @[convert.scala 26:67]
  wire [1:0] _T_206; // @[convert.scala 26:51]
  wire [5:0] _T_207; // @[Cat.scala 29:58]
  wire [4:0] _T_209; // @[convert.scala 29:56]
  wire  _T_210; // @[convert.scala 29:60]
  wire  _T_211; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_214; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [5:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_222; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_223; // @[PositFMA.scala 59:34]
  wire  _T_224; // @[PositFMA.scala 59:47]
  wire  _T_225; // @[PositFMA.scala 59:45]
  wire [2:0] _T_227; // @[Cat.scala 29:58]
  wire [2:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_228; // @[PositFMA.scala 60:34]
  wire  _T_229; // @[PositFMA.scala 60:47]
  wire  _T_230; // @[PositFMA.scala 60:45]
  wire [2:0] _T_232; // @[Cat.scala 29:58]
  wire [2:0] sigB; // @[PositFMA.scala 60:76]
  wire [5:0] _T_233; // @[PositFMA.scala 62:25]
  wire [5:0] sigP; // @[PositFMA.scala 62:33]
  wire [1:0] head2; // @[PositFMA.scala 63:28]
  wire  _T_234; // @[PositFMA.scala 64:31]
  wire  _T_235; // @[PositFMA.scala 64:25]
  wire  _T_236; // @[PositFMA.scala 64:42]
  wire  addTwo; // @[PositFMA.scala 64:35]
  wire  _T_237; // @[PositFMA.scala 66:23]
  wire  _T_238; // @[PositFMA.scala 66:49]
  wire  addOne; // @[PositFMA.scala 66:43]
  wire [1:0] _T_239; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 67:39]
  wire  mulSign; // @[PositFMA.scala 68:28]
  wire [6:0] _T_240; // @[PositFMA.scala 70:30]
  wire [6:0] _GEN_12; // @[PositFMA.scala 70:44]
  wire [6:0] _T_242; // @[PositFMA.scala 70:44]
  wire [6:0] mulScale; // @[PositFMA.scala 70:44]
  wire [3:0] _T_243; // @[PositFMA.scala 73:29]
  wire [2:0] _T_244; // @[PositFMA.scala 74:29]
  wire [3:0] _T_245; // @[PositFMA.scala 74:48]
  wire [3:0] mulSigTmp; // @[PositFMA.scala 71:22]
  wire  _T_247; // @[PositFMA.scala 78:39]
  wire  _T_248; // @[PositFMA.scala 78:43]
  wire [2:0] _T_249; // @[PositFMA.scala 79:39]
  wire [4:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [4:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [6:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [5:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_275; // @[PositFMA.scala 108:29]
  wire  _T_276; // @[PositFMA.scala 108:47]
  wire  _T_277; // @[PositFMA.scala 108:45]
  wire [4:0] extAddSig; // @[Cat.scala 29:58]
  wire [6:0] _GEN_13; // @[PositFMA.scala 112:39]
  wire  mulGreater; // @[PositFMA.scala 112:39]
  wire [6:0] greaterScale; // @[PositFMA.scala 113:26]
  wire [6:0] smallerScale; // @[PositFMA.scala 114:26]
  wire [6:0] _T_281; // @[PositFMA.scala 115:36]
  wire [6:0] scaleDiff; // @[PositFMA.scala 115:36]
  wire [4:0] greaterSig; // @[PositFMA.scala 116:26]
  wire [4:0] smallerSigTmp; // @[PositFMA.scala 117:26]
  wire [6:0] _T_282; // @[PositFMA.scala 118:69]
  wire  _T_283; // @[Shift.scala 39:24]
  wire [2:0] _T_284; // @[Shift.scala 40:44]
  wire  _T_285; // @[Shift.scala 90:30]
  wire [3:0] _T_286; // @[Shift.scala 90:48]
  wire  _T_287; // @[Shift.scala 90:57]
  wire  _T_288; // @[Shift.scala 90:39]
  wire  _T_289; // @[Shift.scala 12:21]
  wire  _T_290; // @[Shift.scala 12:21]
  wire [3:0] _T_292; // @[Bitwise.scala 71:12]
  wire [4:0] _T_293; // @[Cat.scala 29:58]
  wire [4:0] _T_294; // @[Shift.scala 91:22]
  wire [1:0] _T_295; // @[Shift.scala 92:77]
  wire [2:0] _T_296; // @[Shift.scala 90:30]
  wire [1:0] _T_297; // @[Shift.scala 90:48]
  wire  _T_298; // @[Shift.scala 90:57]
  wire [2:0] _GEN_14; // @[Shift.scala 90:39]
  wire [2:0] _T_299; // @[Shift.scala 90:39]
  wire  _T_300; // @[Shift.scala 12:21]
  wire  _T_301; // @[Shift.scala 12:21]
  wire [1:0] _T_303; // @[Bitwise.scala 71:12]
  wire [4:0] _T_304; // @[Cat.scala 29:58]
  wire [4:0] _T_305; // @[Shift.scala 91:22]
  wire  _T_306; // @[Shift.scala 92:77]
  wire [3:0] _T_307; // @[Shift.scala 90:30]
  wire  _T_308; // @[Shift.scala 90:48]
  wire [3:0] _GEN_15; // @[Shift.scala 90:39]
  wire [3:0] _T_310; // @[Shift.scala 90:39]
  wire  _T_312; // @[Shift.scala 12:21]
  wire [4:0] _T_313; // @[Cat.scala 29:58]
  wire [4:0] _T_314; // @[Shift.scala 91:22]
  wire [4:0] _T_317; // @[Bitwise.scala 71:12]
  wire [4:0] smallerSig; // @[Shift.scala 39:10]
  wire [5:0] rawSumSig; // @[PositFMA.scala 119:34]
  wire  _T_318; // @[PositFMA.scala 120:42]
  wire  _T_319; // @[PositFMA.scala 120:46]
  wire  _T_320; // @[PositFMA.scala 120:79]
  wire  sumSign; // @[PositFMA.scala 120:63]
  wire [4:0] _T_322; // @[PositFMA.scala 121:50]
  wire [5:0] signSumSig; // @[Cat.scala 29:58]
  wire [4:0] _T_323; // @[PositFMA.scala 126:33]
  wire [4:0] _T_324; // @[PositFMA.scala 126:68]
  wire [4:0] sumXor; // @[PositFMA.scala 126:51]
  wire [3:0] _T_325; // @[LZD.scala 43:32]
  wire [1:0] _T_326; // @[LZD.scala 43:32]
  wire  _T_327; // @[LZD.scala 39:14]
  wire  _T_328; // @[LZD.scala 39:21]
  wire  _T_329; // @[LZD.scala 39:30]
  wire  _T_330; // @[LZD.scala 39:27]
  wire  _T_331; // @[LZD.scala 39:25]
  wire [1:0] _T_332; // @[Cat.scala 29:58]
  wire [1:0] _T_333; // @[LZD.scala 44:32]
  wire  _T_334; // @[LZD.scala 39:14]
  wire  _T_335; // @[LZD.scala 39:21]
  wire  _T_336; // @[LZD.scala 39:30]
  wire  _T_337; // @[LZD.scala 39:27]
  wire  _T_338; // @[LZD.scala 39:25]
  wire [1:0] _T_339; // @[Cat.scala 29:58]
  wire  _T_340; // @[Shift.scala 12:21]
  wire  _T_341; // @[Shift.scala 12:21]
  wire  _T_342; // @[LZD.scala 49:16]
  wire  _T_343; // @[LZD.scala 49:27]
  wire  _T_344; // @[LZD.scala 49:25]
  wire  _T_345; // @[LZD.scala 49:47]
  wire  _T_346; // @[LZD.scala 49:59]
  wire  _T_347; // @[LZD.scala 49:35]
  wire [2:0] _T_349; // @[Cat.scala 29:58]
  wire  _T_350; // @[LZD.scala 44:32]
  wire  _T_352; // @[Shift.scala 12:21]
  wire [1:0] _T_354; // @[Cat.scala 29:58]
  wire [1:0] _T_355; // @[LZD.scala 55:32]
  wire [1:0] _T_356; // @[LZD.scala 55:20]
  wire [2:0] sumLZD; // @[Cat.scala 29:58]
  wire [2:0] shiftValue; // @[PositFMA.scala 128:24]
  wire [3:0] _T_357; // @[PositFMA.scala 129:38]
  wire  _T_358; // @[Shift.scala 16:24]
  wire [1:0] _T_359; // @[Shift.scala 17:37]
  wire  _T_360; // @[Shift.scala 12:21]
  wire [1:0] _T_361; // @[Shift.scala 64:52]
  wire [3:0] _T_363; // @[Cat.scala 29:58]
  wire [3:0] _T_364; // @[Shift.scala 64:27]
  wire  _T_365; // @[Shift.scala 66:70]
  wire [2:0] _T_367; // @[Shift.scala 64:52]
  wire [3:0] _T_368; // @[Cat.scala 29:58]
  wire [3:0] _T_369; // @[Shift.scala 64:27]
  wire [3:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [6:0] _T_371; // @[PositFMA.scala 132:36]
  wire [6:0] _T_372; // @[PositFMA.scala 132:36]
  wire [3:0] _T_373; // @[Cat.scala 29:58]
  wire [3:0] _T_374; // @[PositFMA.scala 132:61]
  wire [6:0] _GEN_16; // @[PositFMA.scala 132:42]
  wire [6:0] _T_376; // @[PositFMA.scala 132:42]
  wire [6:0] sumScale; // @[PositFMA.scala 132:42]
  wire  sumFrac; // @[PositFMA.scala 133:41]
  wire [2:0] grsTmp; // @[PositFMA.scala 136:41]
  wire [1:0] _T_377; // @[PositFMA.scala 139:40]
  wire  _T_378; // @[PositFMA.scala 139:56]
  wire  underflow; // @[PositFMA.scala 146:32]
  wire  overflow; // @[PositFMA.scala 147:32]
  wire  _T_380; // @[PositFMA.scala 156:32]
  wire  decF_isZero; // @[PositFMA.scala 156:20]
  wire [6:0] _T_382; // @[Mux.scala 87:16]
  wire [6:0] _T_383; // @[Mux.scala 87:16]
  wire [5:0] _GEN_17; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  wire [5:0] decF_scale; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  wire [1:0] _T_384; // @[convert.scala 46:61]
  wire [1:0] _T_385; // @[convert.scala 46:52]
  wire [1:0] _T_387; // @[convert.scala 46:42]
  wire [3:0] _T_388; // @[convert.scala 48:34]
  wire  _T_389; // @[convert.scala 49:36]
  wire [3:0] _T_391; // @[convert.scala 50:36]
  wire [3:0] _T_392; // @[convert.scala 50:36]
  wire [3:0] _T_393; // @[convert.scala 50:28]
  wire  _T_394; // @[convert.scala 51:31]
  wire  _T_395; // @[convert.scala 52:43]
  wire [7:0] _T_399; // @[Cat.scala 29:58]
  wire [3:0] _T_400; // @[Shift.scala 39:17]
  wire  _T_401; // @[Shift.scala 39:24]
  wire [2:0] _T_402; // @[Shift.scala 40:44]
  wire [3:0] _T_403; // @[Shift.scala 90:30]
  wire [3:0] _T_404; // @[Shift.scala 90:48]
  wire  _T_405; // @[Shift.scala 90:57]
  wire [3:0] _GEN_18; // @[Shift.scala 90:39]
  wire [3:0] _T_406; // @[Shift.scala 90:39]
  wire  _T_407; // @[Shift.scala 12:21]
  wire  _T_408; // @[Shift.scala 12:21]
  wire [3:0] _T_410; // @[Bitwise.scala 71:12]
  wire [7:0] _T_411; // @[Cat.scala 29:58]
  wire [7:0] _T_412; // @[Shift.scala 91:22]
  wire [1:0] _T_413; // @[Shift.scala 92:77]
  wire [5:0] _T_414; // @[Shift.scala 90:30]
  wire [1:0] _T_415; // @[Shift.scala 90:48]
  wire  _T_416; // @[Shift.scala 90:57]
  wire [5:0] _GEN_19; // @[Shift.scala 90:39]
  wire [5:0] _T_417; // @[Shift.scala 90:39]
  wire  _T_418; // @[Shift.scala 12:21]
  wire  _T_419; // @[Shift.scala 12:21]
  wire [1:0] _T_421; // @[Bitwise.scala 71:12]
  wire [7:0] _T_422; // @[Cat.scala 29:58]
  wire [7:0] _T_423; // @[Shift.scala 91:22]
  wire  _T_424; // @[Shift.scala 92:77]
  wire [6:0] _T_425; // @[Shift.scala 90:30]
  wire  _T_426; // @[Shift.scala 90:48]
  wire [6:0] _GEN_20; // @[Shift.scala 90:39]
  wire [6:0] _T_428; // @[Shift.scala 90:39]
  wire  _T_430; // @[Shift.scala 12:21]
  wire [7:0] _T_431; // @[Cat.scala 29:58]
  wire [7:0] _T_432; // @[Shift.scala 91:22]
  wire [7:0] _T_435; // @[Bitwise.scala 71:12]
  wire [7:0] _T_436; // @[Shift.scala 39:10]
  wire  _T_437; // @[convert.scala 55:31]
  wire  _T_438; // @[convert.scala 56:31]
  wire  _T_439; // @[convert.scala 57:31]
  wire  _T_440; // @[convert.scala 58:31]
  wire [4:0] _T_441; // @[convert.scala 59:69]
  wire  _T_442; // @[convert.scala 59:81]
  wire  _T_443; // @[convert.scala 59:50]
  wire  _T_445; // @[convert.scala 60:81]
  wire  _T_446; // @[convert.scala 61:44]
  wire  _T_447; // @[convert.scala 61:52]
  wire  _T_448; // @[convert.scala 61:36]
  wire  _T_449; // @[convert.scala 62:63]
  wire  _T_450; // @[convert.scala 62:103]
  wire  _T_451; // @[convert.scala 62:60]
  wire [4:0] _GEN_21; // @[convert.scala 63:56]
  wire [4:0] _T_454; // @[convert.scala 63:56]
  wire [5:0] _T_455; // @[Cat.scala 29:58]
  reg  _T_459; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [5:0] _T_463; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 6'h3f : 6'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{5'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 6'h3f : 6'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{5'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[5]; // @[convert.scala 18:24]
  assign _T_14 = realA[4]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[4:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[3:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[3:2]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19 != 2'h0; // @[LZD.scala 39:14]
  assign _T_21 = _T_19[1]; // @[LZD.scala 39:21]
  assign _T_22 = _T_19[0]; // @[LZD.scala 39:30]
  assign _T_23 = ~ _T_22; // @[LZD.scala 39:27]
  assign _T_24 = _T_21 | _T_23; // @[LZD.scala 39:25]
  assign _T_25 = {_T_20,_T_24}; // @[Cat.scala 29:58]
  assign _T_26 = _T_18[1:0]; // @[LZD.scala 44:32]
  assign _T_27 = _T_26 != 2'h0; // @[LZD.scala 39:14]
  assign _T_28 = _T_26[1]; // @[LZD.scala 39:21]
  assign _T_29 = _T_26[0]; // @[LZD.scala 39:30]
  assign _T_30 = ~ _T_29; // @[LZD.scala 39:27]
  assign _T_31 = _T_28 | _T_30; // @[LZD.scala 39:25]
  assign _T_32 = {_T_27,_T_31}; // @[Cat.scala 29:58]
  assign _T_33 = _T_25[1]; // @[Shift.scala 12:21]
  assign _T_34 = _T_32[1]; // @[Shift.scala 12:21]
  assign _T_35 = _T_33 | _T_34; // @[LZD.scala 49:16]
  assign _T_36 = ~ _T_34; // @[LZD.scala 49:27]
  assign _T_37 = _T_33 | _T_36; // @[LZD.scala 49:25]
  assign _T_38 = _T_25[0:0]; // @[LZD.scala 49:47]
  assign _T_39 = _T_32[0:0]; // @[LZD.scala 49:59]
  assign _T_40 = _T_33 ? _T_38 : _T_39; // @[LZD.scala 49:35]
  assign _T_42 = {_T_35,_T_37,_T_40}; // @[Cat.scala 29:58]
  assign _T_43 = ~ _T_42; // @[convert.scala 21:22]
  assign _T_44 = realA[2:0]; // @[convert.scala 22:36]
  assign _T_45 = _T_43 < 3'h3; // @[Shift.scala 16:24]
  assign _T_46 = _T_43[1:0]; // @[Shift.scala 17:37]
  assign _T_47 = _T_46[1]; // @[Shift.scala 12:21]
  assign _T_48 = _T_44[0:0]; // @[Shift.scala 64:52]
  assign _T_50 = {_T_48,2'h0}; // @[Cat.scala 29:58]
  assign _T_51 = _T_47 ? _T_50 : _T_44; // @[Shift.scala 64:27]
  assign _T_52 = _T_46[0:0]; // @[Shift.scala 66:70]
  assign _T_54 = _T_51[1:0]; // @[Shift.scala 64:52]
  assign _T_55 = {_T_54,1'h0}; // @[Cat.scala 29:58]
  assign _T_56 = _T_52 ? _T_55 : _T_51; // @[Shift.scala 64:27]
  assign _T_57 = _T_45 ? _T_56 : 3'h0; // @[Shift.scala 16:10]
  assign _T_58 = _T_57[2:1]; // @[convert.scala 23:34]
  assign decA_fraction = _T_57[0:0]; // @[convert.scala 24:34]
  assign _T_60 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_62 = _T_15 ? _T_43 : _T_42; // @[convert.scala 25:42]
  assign _T_65 = ~ _T_58; // @[convert.scala 26:67]
  assign _T_66 = _T_13 ? _T_65 : _T_58; // @[convert.scala 26:51]
  assign _T_67 = {_T_60,_T_62,_T_66}; // @[Cat.scala 29:58]
  assign _T_69 = realA[4:0]; // @[convert.scala 29:56]
  assign _T_70 = _T_69 != 5'h0; // @[convert.scala 29:60]
  assign _T_71 = ~ _T_70; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_71; // @[convert.scala 29:39]
  assign _T_74 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_74 & _T_71; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_67); // @[convert.scala 32:24]
  assign _T_83 = io_B[5]; // @[convert.scala 18:24]
  assign _T_84 = io_B[4]; // @[convert.scala 18:40]
  assign _T_85 = _T_83 ^ _T_84; // @[convert.scala 18:36]
  assign _T_86 = io_B[4:1]; // @[convert.scala 19:24]
  assign _T_87 = io_B[3:0]; // @[convert.scala 19:43]
  assign _T_88 = _T_86 ^ _T_87; // @[convert.scala 19:39]
  assign _T_89 = _T_88[3:2]; // @[LZD.scala 43:32]
  assign _T_90 = _T_89 != 2'h0; // @[LZD.scala 39:14]
  assign _T_91 = _T_89[1]; // @[LZD.scala 39:21]
  assign _T_92 = _T_89[0]; // @[LZD.scala 39:30]
  assign _T_93 = ~ _T_92; // @[LZD.scala 39:27]
  assign _T_94 = _T_91 | _T_93; // @[LZD.scala 39:25]
  assign _T_95 = {_T_90,_T_94}; // @[Cat.scala 29:58]
  assign _T_96 = _T_88[1:0]; // @[LZD.scala 44:32]
  assign _T_97 = _T_96 != 2'h0; // @[LZD.scala 39:14]
  assign _T_98 = _T_96[1]; // @[LZD.scala 39:21]
  assign _T_99 = _T_96[0]; // @[LZD.scala 39:30]
  assign _T_100 = ~ _T_99; // @[LZD.scala 39:27]
  assign _T_101 = _T_98 | _T_100; // @[LZD.scala 39:25]
  assign _T_102 = {_T_97,_T_101}; // @[Cat.scala 29:58]
  assign _T_103 = _T_95[1]; // @[Shift.scala 12:21]
  assign _T_104 = _T_102[1]; // @[Shift.scala 12:21]
  assign _T_105 = _T_103 | _T_104; // @[LZD.scala 49:16]
  assign _T_106 = ~ _T_104; // @[LZD.scala 49:27]
  assign _T_107 = _T_103 | _T_106; // @[LZD.scala 49:25]
  assign _T_108 = _T_95[0:0]; // @[LZD.scala 49:47]
  assign _T_109 = _T_102[0:0]; // @[LZD.scala 49:59]
  assign _T_110 = _T_103 ? _T_108 : _T_109; // @[LZD.scala 49:35]
  assign _T_112 = {_T_105,_T_107,_T_110}; // @[Cat.scala 29:58]
  assign _T_113 = ~ _T_112; // @[convert.scala 21:22]
  assign _T_114 = io_B[2:0]; // @[convert.scala 22:36]
  assign _T_115 = _T_113 < 3'h3; // @[Shift.scala 16:24]
  assign _T_116 = _T_113[1:0]; // @[Shift.scala 17:37]
  assign _T_117 = _T_116[1]; // @[Shift.scala 12:21]
  assign _T_118 = _T_114[0:0]; // @[Shift.scala 64:52]
  assign _T_120 = {_T_118,2'h0}; // @[Cat.scala 29:58]
  assign _T_121 = _T_117 ? _T_120 : _T_114; // @[Shift.scala 64:27]
  assign _T_122 = _T_116[0:0]; // @[Shift.scala 66:70]
  assign _T_124 = _T_121[1:0]; // @[Shift.scala 64:52]
  assign _T_125 = {_T_124,1'h0}; // @[Cat.scala 29:58]
  assign _T_126 = _T_122 ? _T_125 : _T_121; // @[Shift.scala 64:27]
  assign _T_127 = _T_115 ? _T_126 : 3'h0; // @[Shift.scala 16:10]
  assign _T_128 = _T_127[2:1]; // @[convert.scala 23:34]
  assign decB_fraction = _T_127[0:0]; // @[convert.scala 24:34]
  assign _T_130 = _T_85 == 1'h0; // @[convert.scala 25:26]
  assign _T_132 = _T_85 ? _T_113 : _T_112; // @[convert.scala 25:42]
  assign _T_135 = ~ _T_128; // @[convert.scala 26:67]
  assign _T_136 = _T_83 ? _T_135 : _T_128; // @[convert.scala 26:51]
  assign _T_137 = {_T_130,_T_132,_T_136}; // @[Cat.scala 29:58]
  assign _T_139 = io_B[4:0]; // @[convert.scala 29:56]
  assign _T_140 = _T_139 != 5'h0; // @[convert.scala 29:60]
  assign _T_141 = ~ _T_140; // @[convert.scala 29:41]
  assign decB_isNaR = _T_83 & _T_141; // @[convert.scala 29:39]
  assign _T_144 = _T_83 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_144 & _T_141; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_137); // @[convert.scala 32:24]
  assign _T_153 = realC[5]; // @[convert.scala 18:24]
  assign _T_154 = realC[4]; // @[convert.scala 18:40]
  assign _T_155 = _T_153 ^ _T_154; // @[convert.scala 18:36]
  assign _T_156 = realC[4:1]; // @[convert.scala 19:24]
  assign _T_157 = realC[3:0]; // @[convert.scala 19:43]
  assign _T_158 = _T_156 ^ _T_157; // @[convert.scala 19:39]
  assign _T_159 = _T_158[3:2]; // @[LZD.scala 43:32]
  assign _T_160 = _T_159 != 2'h0; // @[LZD.scala 39:14]
  assign _T_161 = _T_159[1]; // @[LZD.scala 39:21]
  assign _T_162 = _T_159[0]; // @[LZD.scala 39:30]
  assign _T_163 = ~ _T_162; // @[LZD.scala 39:27]
  assign _T_164 = _T_161 | _T_163; // @[LZD.scala 39:25]
  assign _T_165 = {_T_160,_T_164}; // @[Cat.scala 29:58]
  assign _T_166 = _T_158[1:0]; // @[LZD.scala 44:32]
  assign _T_167 = _T_166 != 2'h0; // @[LZD.scala 39:14]
  assign _T_168 = _T_166[1]; // @[LZD.scala 39:21]
  assign _T_169 = _T_166[0]; // @[LZD.scala 39:30]
  assign _T_170 = ~ _T_169; // @[LZD.scala 39:27]
  assign _T_171 = _T_168 | _T_170; // @[LZD.scala 39:25]
  assign _T_172 = {_T_167,_T_171}; // @[Cat.scala 29:58]
  assign _T_173 = _T_165[1]; // @[Shift.scala 12:21]
  assign _T_174 = _T_172[1]; // @[Shift.scala 12:21]
  assign _T_175 = _T_173 | _T_174; // @[LZD.scala 49:16]
  assign _T_176 = ~ _T_174; // @[LZD.scala 49:27]
  assign _T_177 = _T_173 | _T_176; // @[LZD.scala 49:25]
  assign _T_178 = _T_165[0:0]; // @[LZD.scala 49:47]
  assign _T_179 = _T_172[0:0]; // @[LZD.scala 49:59]
  assign _T_180 = _T_173 ? _T_178 : _T_179; // @[LZD.scala 49:35]
  assign _T_182 = {_T_175,_T_177,_T_180}; // @[Cat.scala 29:58]
  assign _T_183 = ~ _T_182; // @[convert.scala 21:22]
  assign _T_184 = realC[2:0]; // @[convert.scala 22:36]
  assign _T_185 = _T_183 < 3'h3; // @[Shift.scala 16:24]
  assign _T_186 = _T_183[1:0]; // @[Shift.scala 17:37]
  assign _T_187 = _T_186[1]; // @[Shift.scala 12:21]
  assign _T_188 = _T_184[0:0]; // @[Shift.scala 64:52]
  assign _T_190 = {_T_188,2'h0}; // @[Cat.scala 29:58]
  assign _T_191 = _T_187 ? _T_190 : _T_184; // @[Shift.scala 64:27]
  assign _T_192 = _T_186[0:0]; // @[Shift.scala 66:70]
  assign _T_194 = _T_191[1:0]; // @[Shift.scala 64:52]
  assign _T_195 = {_T_194,1'h0}; // @[Cat.scala 29:58]
  assign _T_196 = _T_192 ? _T_195 : _T_191; // @[Shift.scala 64:27]
  assign _T_197 = _T_185 ? _T_196 : 3'h0; // @[Shift.scala 16:10]
  assign _T_198 = _T_197[2:1]; // @[convert.scala 23:34]
  assign decC_fraction = _T_197[0:0]; // @[convert.scala 24:34]
  assign _T_200 = _T_155 == 1'h0; // @[convert.scala 25:26]
  assign _T_202 = _T_155 ? _T_183 : _T_182; // @[convert.scala 25:42]
  assign _T_205 = ~ _T_198; // @[convert.scala 26:67]
  assign _T_206 = _T_153 ? _T_205 : _T_198; // @[convert.scala 26:51]
  assign _T_207 = {_T_200,_T_202,_T_206}; // @[Cat.scala 29:58]
  assign _T_209 = realC[4:0]; // @[convert.scala 29:56]
  assign _T_210 = _T_209 != 5'h0; // @[convert.scala 29:60]
  assign _T_211 = ~ _T_210; // @[convert.scala 29:41]
  assign decC_isNaR = _T_153 & _T_211; // @[convert.scala 29:39]
  assign _T_214 = _T_153 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_214 & _T_211; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_207); // @[convert.scala 32:24]
  assign _T_222 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_222 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_223 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_224 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_225 = _T_223 & _T_224; // @[PositFMA.scala 59:45]
  assign _T_227 = {_T_13,_T_225,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_227); // @[PositFMA.scala 59:76]
  assign _T_228 = ~ _T_83; // @[PositFMA.scala 60:34]
  assign _T_229 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_230 = _T_228 & _T_229; // @[PositFMA.scala 60:45]
  assign _T_232 = {_T_83,_T_230,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_232); // @[PositFMA.scala 60:76]
  assign _T_233 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 62:25]
  assign sigP = $unsigned(_T_233); // @[PositFMA.scala 62:33]
  assign head2 = sigP[5:4]; // @[PositFMA.scala 63:28]
  assign _T_234 = head2[1]; // @[PositFMA.scala 64:31]
  assign _T_235 = ~ _T_234; // @[PositFMA.scala 64:25]
  assign _T_236 = head2[0]; // @[PositFMA.scala 64:42]
  assign addTwo = _T_235 & _T_236; // @[PositFMA.scala 64:35]
  assign _T_237 = sigP[5]; // @[PositFMA.scala 66:23]
  assign _T_238 = sigP[3]; // @[PositFMA.scala 66:49]
  assign addOne = _T_237 ^ _T_238; // @[PositFMA.scala 66:43]
  assign _T_239 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_239)}; // @[PositFMA.scala 67:39]
  assign mulSign = sigP[5:5]; // @[PositFMA.scala 68:28]
  assign _T_240 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 70:30]
  assign _GEN_12 = {{4{expBias[2]}},expBias}; // @[PositFMA.scala 70:44]
  assign _T_242 = $signed(_T_240) + $signed(_GEN_12); // @[PositFMA.scala 70:44]
  assign mulScale = $signed(_T_242); // @[PositFMA.scala 70:44]
  assign _T_243 = sigP[3:0]; // @[PositFMA.scala 73:29]
  assign _T_244 = sigP[2:0]; // @[PositFMA.scala 74:29]
  assign _T_245 = {_T_244, 1'h0}; // @[PositFMA.scala 74:48]
  assign mulSigTmp = addOne ? _T_243 : _T_245; // @[PositFMA.scala 71:22]
  assign _T_247 = mulSigTmp[3:3]; // @[PositFMA.scala 78:39]
  assign _T_248 = _T_247 | addTwo; // @[PositFMA.scala 78:43]
  assign _T_249 = mulSigTmp[2:0]; // @[PositFMA.scala 79:39]
  assign mulSig = {mulSign,_T_248,_T_249}; // @[Cat.scala 29:58]
  assign _T_275 = ~ addSign_phase2; // @[PositFMA.scala 108:29]
  assign _T_276 = ~ addZero_phase2; // @[PositFMA.scala 108:47]
  assign _T_277 = _T_275 & _T_276; // @[PositFMA.scala 108:45]
  assign extAddSig = {addSign_phase2,_T_277,addFrac_phase2,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[5]}},addScale_phase2}; // @[PositFMA.scala 112:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 112:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[5]}},addScale_phase2}); // @[PositFMA.scala 113:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[5]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 114:26]
  assign _T_281 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 115:36]
  assign scaleDiff = $signed(_T_281); // @[PositFMA.scala 115:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 116:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 117:26]
  assign _T_282 = $unsigned(scaleDiff); // @[PositFMA.scala 118:69]
  assign _T_283 = _T_282 < 7'h5; // @[Shift.scala 39:24]
  assign _T_284 = _T_282[2:0]; // @[Shift.scala 40:44]
  assign _T_285 = smallerSigTmp[4:4]; // @[Shift.scala 90:30]
  assign _T_286 = smallerSigTmp[3:0]; // @[Shift.scala 90:48]
  assign _T_287 = _T_286 != 4'h0; // @[Shift.scala 90:57]
  assign _T_288 = _T_285 | _T_287; // @[Shift.scala 90:39]
  assign _T_289 = _T_284[2]; // @[Shift.scala 12:21]
  assign _T_290 = smallerSigTmp[4]; // @[Shift.scala 12:21]
  assign _T_292 = _T_290 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_293 = {_T_292,_T_288}; // @[Cat.scala 29:58]
  assign _T_294 = _T_289 ? _T_293 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_295 = _T_284[1:0]; // @[Shift.scala 92:77]
  assign _T_296 = _T_294[4:2]; // @[Shift.scala 90:30]
  assign _T_297 = _T_294[1:0]; // @[Shift.scala 90:48]
  assign _T_298 = _T_297 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{2'd0}, _T_298}; // @[Shift.scala 90:39]
  assign _T_299 = _T_296 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_300 = _T_295[1]; // @[Shift.scala 12:21]
  assign _T_301 = _T_294[4]; // @[Shift.scala 12:21]
  assign _T_303 = _T_301 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_304 = {_T_303,_T_299}; // @[Cat.scala 29:58]
  assign _T_305 = _T_300 ? _T_304 : _T_294; // @[Shift.scala 91:22]
  assign _T_306 = _T_295[0:0]; // @[Shift.scala 92:77]
  assign _T_307 = _T_305[4:1]; // @[Shift.scala 90:30]
  assign _T_308 = _T_305[0:0]; // @[Shift.scala 90:48]
  assign _GEN_15 = {{3'd0}, _T_308}; // @[Shift.scala 90:39]
  assign _T_310 = _T_307 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_312 = _T_305[4]; // @[Shift.scala 12:21]
  assign _T_313 = {_T_312,_T_310}; // @[Cat.scala 29:58]
  assign _T_314 = _T_306 ? _T_313 : _T_305; // @[Shift.scala 91:22]
  assign _T_317 = _T_290 ? 5'h1f : 5'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_283 ? _T_314 : _T_317; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 119:34]
  assign _T_318 = mulSig_phase2[4:4]; // @[PositFMA.scala 120:42]
  assign _T_319 = _T_318 ^ addSign_phase2; // @[PositFMA.scala 120:46]
  assign _T_320 = rawSumSig[5:5]; // @[PositFMA.scala 120:79]
  assign sumSign = _T_319 ^ _T_320; // @[PositFMA.scala 120:63]
  assign _T_322 = greaterSig + smallerSig; // @[PositFMA.scala 121:50]
  assign signSumSig = {sumSign,_T_322}; // @[Cat.scala 29:58]
  assign _T_323 = signSumSig[5:1]; // @[PositFMA.scala 126:33]
  assign _T_324 = signSumSig[4:0]; // @[PositFMA.scala 126:68]
  assign sumXor = _T_323 ^ _T_324; // @[PositFMA.scala 126:51]
  assign _T_325 = sumXor[4:1]; // @[LZD.scala 43:32]
  assign _T_326 = _T_325[3:2]; // @[LZD.scala 43:32]
  assign _T_327 = _T_326 != 2'h0; // @[LZD.scala 39:14]
  assign _T_328 = _T_326[1]; // @[LZD.scala 39:21]
  assign _T_329 = _T_326[0]; // @[LZD.scala 39:30]
  assign _T_330 = ~ _T_329; // @[LZD.scala 39:27]
  assign _T_331 = _T_328 | _T_330; // @[LZD.scala 39:25]
  assign _T_332 = {_T_327,_T_331}; // @[Cat.scala 29:58]
  assign _T_333 = _T_325[1:0]; // @[LZD.scala 44:32]
  assign _T_334 = _T_333 != 2'h0; // @[LZD.scala 39:14]
  assign _T_335 = _T_333[1]; // @[LZD.scala 39:21]
  assign _T_336 = _T_333[0]; // @[LZD.scala 39:30]
  assign _T_337 = ~ _T_336; // @[LZD.scala 39:27]
  assign _T_338 = _T_335 | _T_337; // @[LZD.scala 39:25]
  assign _T_339 = {_T_334,_T_338}; // @[Cat.scala 29:58]
  assign _T_340 = _T_332[1]; // @[Shift.scala 12:21]
  assign _T_341 = _T_339[1]; // @[Shift.scala 12:21]
  assign _T_342 = _T_340 | _T_341; // @[LZD.scala 49:16]
  assign _T_343 = ~ _T_341; // @[LZD.scala 49:27]
  assign _T_344 = _T_340 | _T_343; // @[LZD.scala 49:25]
  assign _T_345 = _T_332[0:0]; // @[LZD.scala 49:47]
  assign _T_346 = _T_339[0:0]; // @[LZD.scala 49:59]
  assign _T_347 = _T_340 ? _T_345 : _T_346; // @[LZD.scala 49:35]
  assign _T_349 = {_T_342,_T_344,_T_347}; // @[Cat.scala 29:58]
  assign _T_350 = sumXor[0:0]; // @[LZD.scala 44:32]
  assign _T_352 = _T_349[2]; // @[Shift.scala 12:21]
  assign _T_354 = {1'h1,_T_350}; // @[Cat.scala 29:58]
  assign _T_355 = _T_349[1:0]; // @[LZD.scala 55:32]
  assign _T_356 = _T_352 ? _T_355 : _T_354; // @[LZD.scala 55:20]
  assign sumLZD = {_T_352,_T_356}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 128:24]
  assign _T_357 = signSumSig[3:0]; // @[PositFMA.scala 129:38]
  assign _T_358 = shiftValue < 3'h4; // @[Shift.scala 16:24]
  assign _T_359 = shiftValue[1:0]; // @[Shift.scala 17:37]
  assign _T_360 = _T_359[1]; // @[Shift.scala 12:21]
  assign _T_361 = _T_357[1:0]; // @[Shift.scala 64:52]
  assign _T_363 = {_T_361,2'h0}; // @[Cat.scala 29:58]
  assign _T_364 = _T_360 ? _T_363 : _T_357; // @[Shift.scala 64:27]
  assign _T_365 = _T_359[0:0]; // @[Shift.scala 66:70]
  assign _T_367 = _T_364[2:0]; // @[Shift.scala 64:52]
  assign _T_368 = {_T_367,1'h0}; // @[Cat.scala 29:58]
  assign _T_369 = _T_365 ? _T_368 : _T_364; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_358 ? _T_369 : 4'h0; // @[Shift.scala 16:10]
  assign _T_371 = $signed(greaterScale) + $signed(7'sh2); // @[PositFMA.scala 132:36]
  assign _T_372 = $signed(_T_371); // @[PositFMA.scala 132:36]
  assign _T_373 = {1'h1,_T_352,_T_356}; // @[Cat.scala 29:58]
  assign _T_374 = $signed(_T_373); // @[PositFMA.scala 132:61]
  assign _GEN_16 = {{3{_T_374[3]}},_T_374}; // @[PositFMA.scala 132:42]
  assign _T_376 = $signed(_T_372) + $signed(_GEN_16); // @[PositFMA.scala 132:42]
  assign sumScale = $signed(_T_376); // @[PositFMA.scala 132:42]
  assign sumFrac = normalFracTmp[3:3]; // @[PositFMA.scala 133:41]
  assign grsTmp = normalFracTmp[2:0]; // @[PositFMA.scala 136:41]
  assign _T_377 = grsTmp[2:1]; // @[PositFMA.scala 139:40]
  assign _T_378 = grsTmp[0:0]; // @[PositFMA.scala 139:56]
  assign underflow = $signed(sumScale) < $signed(-7'sh11); // @[PositFMA.scala 146:32]
  assign overflow = $signed(sumScale) > $signed(7'sh10); // @[PositFMA.scala 147:32]
  assign _T_380 = signSumSig != 6'h0; // @[PositFMA.scala 156:32]
  assign decF_isZero = ~ _T_380; // @[PositFMA.scala 156:20]
  assign _T_382 = underflow ? $signed(-7'sh11) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_383 = overflow ? $signed(7'sh10) : $signed(_T_382); // @[Mux.scala 87:16]
  assign _GEN_17 = _T_383[5:0]; // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  assign decF_scale = $signed(_GEN_17); // @[PositFMA.scala 153:18 PositFMA.scala 159:17]
  assign _T_384 = decF_scale[1:0]; // @[convert.scala 46:61]
  assign _T_385 = ~ _T_384; // @[convert.scala 46:52]
  assign _T_387 = sumSign ? _T_385 : _T_384; // @[convert.scala 46:42]
  assign _T_388 = decF_scale[5:2]; // @[convert.scala 48:34]
  assign _T_389 = _T_388[3:3]; // @[convert.scala 49:36]
  assign _T_391 = ~ _T_388; // @[convert.scala 50:36]
  assign _T_392 = $signed(_T_391); // @[convert.scala 50:36]
  assign _T_393 = _T_389 ? $signed(_T_392) : $signed(_T_388); // @[convert.scala 50:28]
  assign _T_394 = _T_389 ^ sumSign; // @[convert.scala 51:31]
  assign _T_395 = ~ _T_394; // @[convert.scala 52:43]
  assign _T_399 = {_T_395,_T_394,_T_387,sumFrac,_T_377,_T_378}; // @[Cat.scala 29:58]
  assign _T_400 = $unsigned(_T_393); // @[Shift.scala 39:17]
  assign _T_401 = _T_400 < 4'h8; // @[Shift.scala 39:24]
  assign _T_402 = _T_393[2:0]; // @[Shift.scala 40:44]
  assign _T_403 = _T_399[7:4]; // @[Shift.scala 90:30]
  assign _T_404 = _T_399[3:0]; // @[Shift.scala 90:48]
  assign _T_405 = _T_404 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_18 = {{3'd0}, _T_405}; // @[Shift.scala 90:39]
  assign _T_406 = _T_403 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_407 = _T_402[2]; // @[Shift.scala 12:21]
  assign _T_408 = _T_399[7]; // @[Shift.scala 12:21]
  assign _T_410 = _T_408 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_411 = {_T_410,_T_406}; // @[Cat.scala 29:58]
  assign _T_412 = _T_407 ? _T_411 : _T_399; // @[Shift.scala 91:22]
  assign _T_413 = _T_402[1:0]; // @[Shift.scala 92:77]
  assign _T_414 = _T_412[7:2]; // @[Shift.scala 90:30]
  assign _T_415 = _T_412[1:0]; // @[Shift.scala 90:48]
  assign _T_416 = _T_415 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_19 = {{5'd0}, _T_416}; // @[Shift.scala 90:39]
  assign _T_417 = _T_414 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_418 = _T_413[1]; // @[Shift.scala 12:21]
  assign _T_419 = _T_412[7]; // @[Shift.scala 12:21]
  assign _T_421 = _T_419 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_422 = {_T_421,_T_417}; // @[Cat.scala 29:58]
  assign _T_423 = _T_418 ? _T_422 : _T_412; // @[Shift.scala 91:22]
  assign _T_424 = _T_413[0:0]; // @[Shift.scala 92:77]
  assign _T_425 = _T_423[7:1]; // @[Shift.scala 90:30]
  assign _T_426 = _T_423[0:0]; // @[Shift.scala 90:48]
  assign _GEN_20 = {{6'd0}, _T_426}; // @[Shift.scala 90:39]
  assign _T_428 = _T_425 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_430 = _T_423[7]; // @[Shift.scala 12:21]
  assign _T_431 = {_T_430,_T_428}; // @[Cat.scala 29:58]
  assign _T_432 = _T_424 ? _T_431 : _T_423; // @[Shift.scala 91:22]
  assign _T_435 = _T_408 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_436 = _T_401 ? _T_432 : _T_435; // @[Shift.scala 39:10]
  assign _T_437 = _T_436[3]; // @[convert.scala 55:31]
  assign _T_438 = _T_436[2]; // @[convert.scala 56:31]
  assign _T_439 = _T_436[1]; // @[convert.scala 57:31]
  assign _T_440 = _T_436[0]; // @[convert.scala 58:31]
  assign _T_441 = _T_436[7:3]; // @[convert.scala 59:69]
  assign _T_442 = _T_441 != 5'h0; // @[convert.scala 59:81]
  assign _T_443 = ~ _T_442; // @[convert.scala 59:50]
  assign _T_445 = _T_441 == 5'h1f; // @[convert.scala 60:81]
  assign _T_446 = _T_437 | _T_439; // @[convert.scala 61:44]
  assign _T_447 = _T_446 | _T_440; // @[convert.scala 61:52]
  assign _T_448 = _T_438 & _T_447; // @[convert.scala 61:36]
  assign _T_449 = ~ _T_445; // @[convert.scala 62:63]
  assign _T_450 = _T_449 & _T_448; // @[convert.scala 62:103]
  assign _T_451 = _T_443 | _T_450; // @[convert.scala 62:60]
  assign _GEN_21 = {{4'd0}, _T_451}; // @[convert.scala 63:56]
  assign _T_454 = _T_441 + _GEN_21; // @[convert.scala 63:56]
  assign _T_455 = {sumSign,_T_454}; // @[Cat.scala 29:58]
  assign io_F = _T_463; // @[PositFMA.scala 176:15]
  assign io_outValid = _T_459; // @[PositFMA.scala 175:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulSig_phase2 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_459 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_463 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_153;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_459 <= 1'h0;
    end else begin
      _T_459 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_463 <= 6'h20;
      end else begin
        if (decF_isZero) begin
          _T_463 <= 6'h0;
        end else begin
          _T_463 <= _T_455;
        end
      end
    end
  end
endmodule
