module PositMulDec6_0(
  input        clock,
  input        reset,
  input  [5:0] io_A,
  input  [5:0] io_B,
  output [4:0] io_sigA,
  output [4:0] io_sigB,
  output [3:0] io_decAscale,
  output [3:0] io_decBscale,
  output       io_decAisNar,
  output       io_decBisNar,
  output       io_decAisZero,
  output       io_decBisZero
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [3:0] _T_4; // @[convert.scala 19:24]
  wire [3:0] _T_5; // @[convert.scala 19:43]
  wire [3:0] _T_6; // @[convert.scala 19:39]
  wire [1:0] _T_7; // @[LZD.scala 43:32]
  wire  _T_8; // @[LZD.scala 39:14]
  wire  _T_9; // @[LZD.scala 39:21]
  wire  _T_10; // @[LZD.scala 39:30]
  wire  _T_11; // @[LZD.scala 39:27]
  wire  _T_12; // @[LZD.scala 39:25]
  wire [1:0] _T_13; // @[Cat.scala 29:58]
  wire [1:0] _T_14; // @[LZD.scala 44:32]
  wire  _T_15; // @[LZD.scala 39:14]
  wire  _T_16; // @[LZD.scala 39:21]
  wire  _T_17; // @[LZD.scala 39:30]
  wire  _T_18; // @[LZD.scala 39:27]
  wire  _T_19; // @[LZD.scala 39:25]
  wire [1:0] _T_20; // @[Cat.scala 29:58]
  wire  _T_21; // @[Shift.scala 12:21]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[LZD.scala 49:16]
  wire  _T_24; // @[LZD.scala 49:27]
  wire  _T_25; // @[LZD.scala 49:25]
  wire  _T_26; // @[LZD.scala 49:47]
  wire  _T_27; // @[LZD.scala 49:59]
  wire  _T_28; // @[LZD.scala 49:35]
  wire [2:0] _T_30; // @[Cat.scala 29:58]
  wire [2:0] _T_31; // @[convert.scala 21:22]
  wire [2:0] _T_32; // @[convert.scala 22:36]
  wire  _T_33; // @[Shift.scala 16:24]
  wire [1:0] _T_34; // @[Shift.scala 17:37]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[Shift.scala 64:52]
  wire [2:0] _T_38; // @[Cat.scala 29:58]
  wire [2:0] _T_39; // @[Shift.scala 64:27]
  wire  _T_40; // @[Shift.scala 66:70]
  wire [1:0] _T_42; // @[Shift.scala 64:52]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire [2:0] _T_44; // @[Shift.scala 64:27]
  wire [2:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_48; // @[convert.scala 25:26]
  wire [2:0] _T_50; // @[convert.scala 25:42]
  wire [3:0] _T_51; // @[Cat.scala 29:58]
  wire [4:0] _T_53; // @[convert.scala 29:56]
  wire  _T_54; // @[convert.scala 29:60]
  wire  _T_55; // @[convert.scala 29:41]
  wire  _T_58; // @[convert.scala 30:19]
  wire  _T_67; // @[convert.scala 18:24]
  wire  _T_68; // @[convert.scala 18:40]
  wire  _T_69; // @[convert.scala 18:36]
  wire [3:0] _T_70; // @[convert.scala 19:24]
  wire [3:0] _T_71; // @[convert.scala 19:43]
  wire [3:0] _T_72; // @[convert.scala 19:39]
  wire [1:0] _T_73; // @[LZD.scala 43:32]
  wire  _T_74; // @[LZD.scala 39:14]
  wire  _T_75; // @[LZD.scala 39:21]
  wire  _T_76; // @[LZD.scala 39:30]
  wire  _T_77; // @[LZD.scala 39:27]
  wire  _T_78; // @[LZD.scala 39:25]
  wire [1:0] _T_79; // @[Cat.scala 29:58]
  wire [1:0] _T_80; // @[LZD.scala 44:32]
  wire  _T_81; // @[LZD.scala 39:14]
  wire  _T_82; // @[LZD.scala 39:21]
  wire  _T_83; // @[LZD.scala 39:30]
  wire  _T_84; // @[LZD.scala 39:27]
  wire  _T_85; // @[LZD.scala 39:25]
  wire [1:0] _T_86; // @[Cat.scala 29:58]
  wire  _T_87; // @[Shift.scala 12:21]
  wire  _T_88; // @[Shift.scala 12:21]
  wire  _T_89; // @[LZD.scala 49:16]
  wire  _T_90; // @[LZD.scala 49:27]
  wire  _T_91; // @[LZD.scala 49:25]
  wire  _T_92; // @[LZD.scala 49:47]
  wire  _T_93; // @[LZD.scala 49:59]
  wire  _T_94; // @[LZD.scala 49:35]
  wire [2:0] _T_96; // @[Cat.scala 29:58]
  wire [2:0] _T_97; // @[convert.scala 21:22]
  wire [2:0] _T_98; // @[convert.scala 22:36]
  wire  _T_99; // @[Shift.scala 16:24]
  wire [1:0] _T_100; // @[Shift.scala 17:37]
  wire  _T_101; // @[Shift.scala 12:21]
  wire  _T_102; // @[Shift.scala 64:52]
  wire [2:0] _T_104; // @[Cat.scala 29:58]
  wire [2:0] _T_105; // @[Shift.scala 64:27]
  wire  _T_106; // @[Shift.scala 66:70]
  wire [1:0] _T_108; // @[Shift.scala 64:52]
  wire [2:0] _T_109; // @[Cat.scala 29:58]
  wire [2:0] _T_110; // @[Shift.scala 64:27]
  wire [2:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_114; // @[convert.scala 25:26]
  wire [2:0] _T_116; // @[convert.scala 25:42]
  wire [3:0] _T_117; // @[Cat.scala 29:58]
  wire [4:0] _T_119; // @[convert.scala 29:56]
  wire  _T_120; // @[convert.scala 29:60]
  wire  _T_121; // @[convert.scala 29:41]
  wire  _T_124; // @[convert.scala 30:19]
  wire  _T_132; // @[PositMulDec.scala 31:34]
  wire [4:0] _T_134; // @[Cat.scala 29:58]
  wire  _T_136; // @[PositMulDec.scala 32:34]
  wire [4:0] _T_138; // @[Cat.scala 29:58]
  assign _T_1 = io_A[5]; // @[convert.scala 18:24]
  assign _T_2 = io_A[4]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[4:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[3:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[3:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7 != 2'h0; // @[LZD.scala 39:14]
  assign _T_9 = _T_7[1]; // @[LZD.scala 39:21]
  assign _T_10 = _T_7[0]; // @[LZD.scala 39:30]
  assign _T_11 = ~ _T_10; // @[LZD.scala 39:27]
  assign _T_12 = _T_9 | _T_11; // @[LZD.scala 39:25]
  assign _T_13 = {_T_8,_T_12}; // @[Cat.scala 29:58]
  assign _T_14 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_15 = _T_14 != 2'h0; // @[LZD.scala 39:14]
  assign _T_16 = _T_14[1]; // @[LZD.scala 39:21]
  assign _T_17 = _T_14[0]; // @[LZD.scala 39:30]
  assign _T_18 = ~ _T_17; // @[LZD.scala 39:27]
  assign _T_19 = _T_16 | _T_18; // @[LZD.scala 39:25]
  assign _T_20 = {_T_15,_T_19}; // @[Cat.scala 29:58]
  assign _T_21 = _T_13[1]; // @[Shift.scala 12:21]
  assign _T_22 = _T_20[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21 | _T_22; // @[LZD.scala 49:16]
  assign _T_24 = ~ _T_22; // @[LZD.scala 49:27]
  assign _T_25 = _T_21 | _T_24; // @[LZD.scala 49:25]
  assign _T_26 = _T_13[0:0]; // @[LZD.scala 49:47]
  assign _T_27 = _T_20[0:0]; // @[LZD.scala 49:59]
  assign _T_28 = _T_21 ? _T_26 : _T_27; // @[LZD.scala 49:35]
  assign _T_30 = {_T_23,_T_25,_T_28}; // @[Cat.scala 29:58]
  assign _T_31 = ~ _T_30; // @[convert.scala 21:22]
  assign _T_32 = io_A[2:0]; // @[convert.scala 22:36]
  assign _T_33 = _T_31 < 3'h3; // @[Shift.scala 16:24]
  assign _T_34 = _T_31[1:0]; // @[Shift.scala 17:37]
  assign _T_35 = _T_34[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_32[0:0]; // @[Shift.scala 64:52]
  assign _T_38 = {_T_36,2'h0}; // @[Cat.scala 29:58]
  assign _T_39 = _T_35 ? _T_38 : _T_32; // @[Shift.scala 64:27]
  assign _T_40 = _T_34[0:0]; // @[Shift.scala 66:70]
  assign _T_42 = _T_39[1:0]; // @[Shift.scala 64:52]
  assign _T_43 = {_T_42,1'h0}; // @[Cat.scala 29:58]
  assign _T_44 = _T_40 ? _T_43 : _T_39; // @[Shift.scala 64:27]
  assign decA_fraction = _T_33 ? _T_44 : 3'h0; // @[Shift.scala 16:10]
  assign _T_48 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_50 = _T_3 ? _T_31 : _T_30; // @[convert.scala 25:42]
  assign _T_51 = {_T_48,_T_50}; // @[Cat.scala 29:58]
  assign _T_53 = io_A[4:0]; // @[convert.scala 29:56]
  assign _T_54 = _T_53 != 5'h0; // @[convert.scala 29:60]
  assign _T_55 = ~ _T_54; // @[convert.scala 29:41]
  assign _T_58 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign _T_67 = io_B[5]; // @[convert.scala 18:24]
  assign _T_68 = io_B[4]; // @[convert.scala 18:40]
  assign _T_69 = _T_67 ^ _T_68; // @[convert.scala 18:36]
  assign _T_70 = io_B[4:1]; // @[convert.scala 19:24]
  assign _T_71 = io_B[3:0]; // @[convert.scala 19:43]
  assign _T_72 = _T_70 ^ _T_71; // @[convert.scala 19:39]
  assign _T_73 = _T_72[3:2]; // @[LZD.scala 43:32]
  assign _T_74 = _T_73 != 2'h0; // @[LZD.scala 39:14]
  assign _T_75 = _T_73[1]; // @[LZD.scala 39:21]
  assign _T_76 = _T_73[0]; // @[LZD.scala 39:30]
  assign _T_77 = ~ _T_76; // @[LZD.scala 39:27]
  assign _T_78 = _T_75 | _T_77; // @[LZD.scala 39:25]
  assign _T_79 = {_T_74,_T_78}; // @[Cat.scala 29:58]
  assign _T_80 = _T_72[1:0]; // @[LZD.scala 44:32]
  assign _T_81 = _T_80 != 2'h0; // @[LZD.scala 39:14]
  assign _T_82 = _T_80[1]; // @[LZD.scala 39:21]
  assign _T_83 = _T_80[0]; // @[LZD.scala 39:30]
  assign _T_84 = ~ _T_83; // @[LZD.scala 39:27]
  assign _T_85 = _T_82 | _T_84; // @[LZD.scala 39:25]
  assign _T_86 = {_T_81,_T_85}; // @[Cat.scala 29:58]
  assign _T_87 = _T_79[1]; // @[Shift.scala 12:21]
  assign _T_88 = _T_86[1]; // @[Shift.scala 12:21]
  assign _T_89 = _T_87 | _T_88; // @[LZD.scala 49:16]
  assign _T_90 = ~ _T_88; // @[LZD.scala 49:27]
  assign _T_91 = _T_87 | _T_90; // @[LZD.scala 49:25]
  assign _T_92 = _T_79[0:0]; // @[LZD.scala 49:47]
  assign _T_93 = _T_86[0:0]; // @[LZD.scala 49:59]
  assign _T_94 = _T_87 ? _T_92 : _T_93; // @[LZD.scala 49:35]
  assign _T_96 = {_T_89,_T_91,_T_94}; // @[Cat.scala 29:58]
  assign _T_97 = ~ _T_96; // @[convert.scala 21:22]
  assign _T_98 = io_B[2:0]; // @[convert.scala 22:36]
  assign _T_99 = _T_97 < 3'h3; // @[Shift.scala 16:24]
  assign _T_100 = _T_97[1:0]; // @[Shift.scala 17:37]
  assign _T_101 = _T_100[1]; // @[Shift.scala 12:21]
  assign _T_102 = _T_98[0:0]; // @[Shift.scala 64:52]
  assign _T_104 = {_T_102,2'h0}; // @[Cat.scala 29:58]
  assign _T_105 = _T_101 ? _T_104 : _T_98; // @[Shift.scala 64:27]
  assign _T_106 = _T_100[0:0]; // @[Shift.scala 66:70]
  assign _T_108 = _T_105[1:0]; // @[Shift.scala 64:52]
  assign _T_109 = {_T_108,1'h0}; // @[Cat.scala 29:58]
  assign _T_110 = _T_106 ? _T_109 : _T_105; // @[Shift.scala 64:27]
  assign decB_fraction = _T_99 ? _T_110 : 3'h0; // @[Shift.scala 16:10]
  assign _T_114 = _T_69 == 1'h0; // @[convert.scala 25:26]
  assign _T_116 = _T_69 ? _T_97 : _T_96; // @[convert.scala 25:42]
  assign _T_117 = {_T_114,_T_116}; // @[Cat.scala 29:58]
  assign _T_119 = io_B[4:0]; // @[convert.scala 29:56]
  assign _T_120 = _T_119 != 5'h0; // @[convert.scala 29:60]
  assign _T_121 = ~ _T_120; // @[convert.scala 29:41]
  assign _T_124 = _T_67 == 1'h0; // @[convert.scala 30:19]
  assign _T_132 = ~ _T_1; // @[PositMulDec.scala 31:34]
  assign _T_134 = {_T_1,_T_132,decA_fraction}; // @[Cat.scala 29:58]
  assign _T_136 = ~ _T_67; // @[PositMulDec.scala 32:34]
  assign _T_138 = {_T_67,_T_136,decB_fraction}; // @[Cat.scala 29:58]
  assign io_sigA = $signed(_T_134); // @[PositMulDec.scala 31:16]
  assign io_sigB = $signed(_T_138); // @[PositMulDec.scala 32:16]
  assign io_decAscale = $signed(_T_51); // @[PositMulDec.scala 33:16]
  assign io_decBscale = $signed(_T_117); // @[PositMulDec.scala 34:16]
  assign io_decAisNar = _T_1 & _T_55; // @[PositMulDec.scala 35:16]
  assign io_decBisNar = _T_67 & _T_121; // @[PositMulDec.scala 36:16]
  assign io_decAisZero = _T_58 & _T_55; // @[PositMulDec.scala 37:17]
  assign io_decBisZero = _T_124 & _T_121; // @[PositMulDec.scala 38:17]
endmodule
