module PositDivSqrter8_4(
  input        clock,
  input        reset,
  output       io_inReady,
  input        io_inValid,
  input        io_sqrtOp,
  input  [7:0] io_A,
  input  [7:0] io_B,
  output       io_diviValid,
  output       io_sqrtValid,
  output       io_invalidExc,
  output [7:0] io_Q
);
  reg [2:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [8:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg  fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [7:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [7:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [5:0] _T_4; // @[convert.scala 19:24]
  wire [5:0] _T_5; // @[convert.scala 19:43]
  wire [5:0] _T_6; // @[convert.scala 19:39]
  wire [3:0] _T_7; // @[LZD.scala 43:32]
  wire [1:0] _T_8; // @[LZD.scala 43:32]
  wire  _T_9; // @[LZD.scala 39:14]
  wire  _T_10; // @[LZD.scala 39:21]
  wire  _T_11; // @[LZD.scala 39:30]
  wire  _T_12; // @[LZD.scala 39:27]
  wire  _T_13; // @[LZD.scala 39:25]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [1:0] _T_15; // @[LZD.scala 44:32]
  wire  _T_16; // @[LZD.scala 39:14]
  wire  _T_17; // @[LZD.scala 39:21]
  wire  _T_18; // @[LZD.scala 39:30]
  wire  _T_19; // @[LZD.scala 39:27]
  wire  _T_20; // @[LZD.scala 39:25]
  wire [1:0] _T_21; // @[Cat.scala 29:58]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[LZD.scala 49:16]
  wire  _T_25; // @[LZD.scala 49:27]
  wire  _T_26; // @[LZD.scala 49:25]
  wire  _T_27; // @[LZD.scala 49:47]
  wire  _T_28; // @[LZD.scala 49:59]
  wire  _T_29; // @[LZD.scala 49:35]
  wire [2:0] _T_31; // @[Cat.scala 29:58]
  wire [1:0] _T_32; // @[LZD.scala 44:32]
  wire  _T_33; // @[LZD.scala 39:14]
  wire  _T_34; // @[LZD.scala 39:21]
  wire  _T_35; // @[LZD.scala 39:30]
  wire  _T_36; // @[LZD.scala 39:27]
  wire  _T_37; // @[LZD.scala 39:25]
  wire [1:0] _T_38; // @[Cat.scala 29:58]
  wire  _T_39; // @[Shift.scala 12:21]
  wire [1:0] _T_41; // @[LZD.scala 55:32]
  wire [1:0] _T_42; // @[LZD.scala 55:20]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire [2:0] _T_44; // @[convert.scala 21:22]
  wire [4:0] _T_45; // @[convert.scala 22:36]
  wire  _T_46; // @[Shift.scala 16:24]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 64:52]
  wire [4:0] _T_51; // @[Cat.scala 29:58]
  wire [4:0] _T_52; // @[Shift.scala 64:27]
  wire [1:0] _T_53; // @[Shift.scala 66:70]
  wire  _T_54; // @[Shift.scala 12:21]
  wire [2:0] _T_55; // @[Shift.scala 64:52]
  wire [4:0] _T_57; // @[Cat.scala 29:58]
  wire [4:0] _T_58; // @[Shift.scala 64:27]
  wire  _T_59; // @[Shift.scala 66:70]
  wire [3:0] _T_61; // @[Shift.scala 64:52]
  wire [4:0] _T_62; // @[Cat.scala 29:58]
  wire [4:0] _T_63; // @[Shift.scala 64:27]
  wire [4:0] _T_64; // @[Shift.scala 16:10]
  wire [3:0] _T_65; // @[convert.scala 23:34]
  wire  decA_fraction; // @[convert.scala 24:34]
  wire  _T_67; // @[convert.scala 25:26]
  wire [2:0] _T_69; // @[convert.scala 25:42]
  wire [3:0] _T_72; // @[convert.scala 26:67]
  wire [3:0] _T_73; // @[convert.scala 26:51]
  wire [7:0] _T_74; // @[Cat.scala 29:58]
  wire [6:0] _T_76; // @[convert.scala 29:56]
  wire  _T_77; // @[convert.scala 29:60]
  wire  _T_78; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_81; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [7:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_90; // @[convert.scala 18:24]
  wire  _T_91; // @[convert.scala 18:40]
  wire  _T_92; // @[convert.scala 18:36]
  wire [5:0] _T_93; // @[convert.scala 19:24]
  wire [5:0] _T_94; // @[convert.scala 19:43]
  wire [5:0] _T_95; // @[convert.scala 19:39]
  wire [3:0] _T_96; // @[LZD.scala 43:32]
  wire [1:0] _T_97; // @[LZD.scala 43:32]
  wire  _T_98; // @[LZD.scala 39:14]
  wire  _T_99; // @[LZD.scala 39:21]
  wire  _T_100; // @[LZD.scala 39:30]
  wire  _T_101; // @[LZD.scala 39:27]
  wire  _T_102; // @[LZD.scala 39:25]
  wire [1:0] _T_103; // @[Cat.scala 29:58]
  wire [1:0] _T_104; // @[LZD.scala 44:32]
  wire  _T_105; // @[LZD.scala 39:14]
  wire  _T_106; // @[LZD.scala 39:21]
  wire  _T_107; // @[LZD.scala 39:30]
  wire  _T_108; // @[LZD.scala 39:27]
  wire  _T_109; // @[LZD.scala 39:25]
  wire [1:0] _T_110; // @[Cat.scala 29:58]
  wire  _T_111; // @[Shift.scala 12:21]
  wire  _T_112; // @[Shift.scala 12:21]
  wire  _T_113; // @[LZD.scala 49:16]
  wire  _T_114; // @[LZD.scala 49:27]
  wire  _T_115; // @[LZD.scala 49:25]
  wire  _T_116; // @[LZD.scala 49:47]
  wire  _T_117; // @[LZD.scala 49:59]
  wire  _T_118; // @[LZD.scala 49:35]
  wire [2:0] _T_120; // @[Cat.scala 29:58]
  wire [1:0] _T_121; // @[LZD.scala 44:32]
  wire  _T_122; // @[LZD.scala 39:14]
  wire  _T_123; // @[LZD.scala 39:21]
  wire  _T_124; // @[LZD.scala 39:30]
  wire  _T_125; // @[LZD.scala 39:27]
  wire  _T_126; // @[LZD.scala 39:25]
  wire [1:0] _T_127; // @[Cat.scala 29:58]
  wire  _T_128; // @[Shift.scala 12:21]
  wire [1:0] _T_130; // @[LZD.scala 55:32]
  wire [1:0] _T_131; // @[LZD.scala 55:20]
  wire [2:0] _T_132; // @[Cat.scala 29:58]
  wire [2:0] _T_133; // @[convert.scala 21:22]
  wire [4:0] _T_134; // @[convert.scala 22:36]
  wire  _T_135; // @[Shift.scala 16:24]
  wire  _T_137; // @[Shift.scala 12:21]
  wire  _T_138; // @[Shift.scala 64:52]
  wire [4:0] _T_140; // @[Cat.scala 29:58]
  wire [4:0] _T_141; // @[Shift.scala 64:27]
  wire [1:0] _T_142; // @[Shift.scala 66:70]
  wire  _T_143; // @[Shift.scala 12:21]
  wire [2:0] _T_144; // @[Shift.scala 64:52]
  wire [4:0] _T_146; // @[Cat.scala 29:58]
  wire [4:0] _T_147; // @[Shift.scala 64:27]
  wire  _T_148; // @[Shift.scala 66:70]
  wire [3:0] _T_150; // @[Shift.scala 64:52]
  wire [4:0] _T_151; // @[Cat.scala 29:58]
  wire [4:0] _T_152; // @[Shift.scala 64:27]
  wire [4:0] _T_153; // @[Shift.scala 16:10]
  wire [3:0] _T_154; // @[convert.scala 23:34]
  wire  decB_fraction; // @[convert.scala 24:34]
  wire  _T_156; // @[convert.scala 25:26]
  wire [2:0] _T_158; // @[convert.scala 25:42]
  wire [3:0] _T_161; // @[convert.scala 26:67]
  wire [3:0] _T_162; // @[convert.scala 26:51]
  wire [7:0] _T_163; // @[Cat.scala 29:58]
  wire [6:0] _T_165; // @[convert.scala 29:56]
  wire  _T_166; // @[convert.scala 29:60]
  wire  _T_167; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_170; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [7:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_179; // @[Bitwise.scala 71:12]
  wire  _T_180; // @[PositDivisionSqrt.scala 80:40]
  wire [7:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_183; // @[PositDivisionSqrt.scala 82:31]
  wire [7:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_186; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_187; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_188; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_189; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_190; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_191; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_192; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_193; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_194; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_195; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [8:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_198; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_199; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_200; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_201; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_202; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_203; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_204; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_205; // @[PositDivisionSqrt.scala 117:30]
  wire [3:0] _T_207; // @[PositDivisionSqrt.scala 119:26]
  wire [3:0] _T_208; // @[PositDivisionSqrt.scala 118:20]
  wire [3:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [3:0] _T_209; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_211; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_212; // @[PositDivisionSqrt.scala 123:27]
  wire [2:0] _T_214; // @[PositDivisionSqrt.scala 123:52]
  wire [2:0] _T_215; // @[PositDivisionSqrt.scala 123:20]
  wire [3:0] _GEN_10; // @[PositDivisionSqrt.scala 122:64]
  wire [3:0] _T_216; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_218; // @[PositDivisionSqrt.scala 124:27]
  wire [3:0] _GEN_11; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _T_220; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _GEN_0; // @[PositDivisionSqrt.scala 116:29]
  wire [6:0] _T_221; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_223; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_224; // @[PositDivisionSqrt.scala 137:28]
  wire [7:0] _T_225; // @[PositDivisionSqrt.scala 146:22]
  wire [5:0] _T_226; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_227; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_228; // @[PositDivisionSqrt.scala 148:23]
  wire [7:0] _T_229; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_230; // @[PositDivisionSqrt.scala 149:23]
  wire [8:0] _T_231; // @[PositDivisionSqrt.scala 149:46]
  wire [7:0] _T_232; // @[PositDivisionSqrt.scala 149:56]
  wire [7:0] _T_233; // @[PositDivisionSqrt.scala 149:16]
  wire [7:0] _T_234; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_235; // @[PositDivisionSqrt.scala 150:17]
  wire [7:0] _T_236; // @[PositDivisionSqrt.scala 150:16]
  wire [7:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_238; // @[PositDivisionSqrt.scala 152:29]
  wire [7:0] _T_239; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_240; // @[PositDivisionSqrt.scala 153:29]
  wire [4:0] _T_241; // @[PositDivisionSqrt.scala 153:22]
  wire [7:0] _GEN_12; // @[PositDivisionSqrt.scala 152:93]
  wire [7:0] _T_242; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_244; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_245; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_246; // @[PositDivisionSqrt.scala 154:57]
  wire [7:0] _T_249; // @[Cat.scala 29:58]
  wire [7:0] _T_250; // @[PositDivisionSqrt.scala 154:22]
  wire [7:0] _T_251; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_253; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_254; // @[PositDivisionSqrt.scala 156:83]
  wire [3:0] _T_256; // @[Bitwise.scala 71:12]
  wire [6:0] bitMask; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  wire [6:0] _GEN_13; // @[PositDivisionSqrt.scala 156:53]
  wire [6:0] _T_257; // @[PositDivisionSqrt.scala 156:53]
  wire [7:0] _GEN_14; // @[PositDivisionSqrt.scala 155:51]
  wire [7:0] _T_258; // @[PositDivisionSqrt.scala 155:51]
  wire [5:0] _T_259; // @[PositDivisionSqrt.scala 157:53]
  wire [7:0] _GEN_15; // @[PositDivisionSqrt.scala 156:89]
  wire [7:0] _T_260; // @[PositDivisionSqrt.scala 156:89]
  wire [7:0] _T_261; // @[PositDivisionSqrt.scala 155:22]
  wire [7:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_263; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_264; // @[PositDivisionSqrt.scala 162:40]
  wire [7:0] _T_267; // @[PositDivisionSqrt.scala 163:97]
  wire [7:0] _T_269; // @[PositDivisionSqrt.scala 164:97]
  wire [7:0] _T_270; // @[PositDivisionSqrt.scala 161:92]
  wire [8:0] _T_275; // @[PositDivisionSqrt.scala 168:98]
  wire [7:0] _T_276; // @[PositDivisionSqrt.scala 168:108]
  wire [7:0] _T_278; // @[PositDivisionSqrt.scala 168:112]
  wire [7:0] _T_282; // @[PositDivisionSqrt.scala 169:112]
  wire [7:0] _T_283; // @[PositDivisionSqrt.scala 166:26]
  wire [7:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_284; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_285; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_287; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_288; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_289; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_290; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_291; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_293; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_294; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_295; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_296; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_297; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_300; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_301; // @[PositDivisionSqrt.scala 187:28]
  wire [7:0] _T_304; // @[PositDivisionSqrt.scala 188:47]
  wire [7:0] _T_305; // @[PositDivisionSqrt.scala 188:18]
  wire [5:0] _T_307; // @[PositDivisionSqrt.scala 189:18]
  wire [7:0] _GEN_16; // @[PositDivisionSqrt.scala 188:78]
  wire [7:0] _T_308; // @[PositDivisionSqrt.scala 188:78]
  wire [7:0] _GEN_17; // @[PositDivisionSqrt.scala 190:47]
  wire [7:0] _T_310; // @[PositDivisionSqrt.scala 190:47]
  wire [7:0] _T_311; // @[PositDivisionSqrt.scala 190:18]
  wire [7:0] _T_312; // @[PositDivisionSqrt.scala 189:78]
  wire [1:0] _T_314; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [7:0] _GEN_18; // @[PositDivisionSqrt.scala 197:25]
  wire [7:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire  _T_317; // @[PositDivisionSqrt.scala 200:97]
  wire  _T_318; // @[PositDivisionSqrt.scala 201:97]
  wire  realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_319; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_320; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_321; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_324; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_325; // @[Cat.scala 29:58]
  wire [2:0] _T_326; // @[PositDivisionSqrt.scala 209:63]
  wire [8:0] _GEN_19; // @[PositDivisionSqrt.scala 209:31]
  wire [8:0] _T_328; // @[PositDivisionSqrt.scala 209:31]
  wire [8:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [8:0] _T_330; // @[Mux.scala 87:16]
  wire [8:0] _T_331; // @[Mux.scala 87:16]
  wire [2:0] _T_332; // @[PositDivisionSqrt.scala 224:48]
  wire [2:0] _T_333; // @[PositDivisionSqrt.scala 224:64]
  wire [2:0] decQ_grs; // @[PositDivisionSqrt.scala 224:23]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [7:0] _GEN_20; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [7:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [3:0] _T_339; // @[convert.scala 46:61]
  wire [3:0] _T_340; // @[convert.scala 46:52]
  wire [3:0] _T_342; // @[convert.scala 46:42]
  wire [3:0] _T_343; // @[convert.scala 48:34]
  wire  _T_344; // @[convert.scala 49:36]
  wire [3:0] _T_346; // @[convert.scala 50:36]
  wire [3:0] _T_347; // @[convert.scala 50:36]
  wire [3:0] _T_348; // @[convert.scala 50:28]
  wire  _T_349; // @[convert.scala 51:31]
  wire  _T_350; // @[convert.scala 52:43]
  wire [9:0] _T_354; // @[Cat.scala 29:58]
  wire [3:0] _T_355; // @[Shift.scala 39:17]
  wire  _T_356; // @[Shift.scala 39:24]
  wire [1:0] _T_358; // @[Shift.scala 90:30]
  wire [7:0] _T_359; // @[Shift.scala 90:48]
  wire  _T_360; // @[Shift.scala 90:57]
  wire [1:0] _GEN_21; // @[Shift.scala 90:39]
  wire [1:0] _T_361; // @[Shift.scala 90:39]
  wire  _T_362; // @[Shift.scala 12:21]
  wire  _T_363; // @[Shift.scala 12:21]
  wire [7:0] _T_365; // @[Bitwise.scala 71:12]
  wire [9:0] _T_366; // @[Cat.scala 29:58]
  wire [9:0] _T_367; // @[Shift.scala 91:22]
  wire [2:0] _T_368; // @[Shift.scala 92:77]
  wire [5:0] _T_369; // @[Shift.scala 90:30]
  wire [3:0] _T_370; // @[Shift.scala 90:48]
  wire  _T_371; // @[Shift.scala 90:57]
  wire [5:0] _GEN_22; // @[Shift.scala 90:39]
  wire [5:0] _T_372; // @[Shift.scala 90:39]
  wire  _T_373; // @[Shift.scala 12:21]
  wire  _T_374; // @[Shift.scala 12:21]
  wire [3:0] _T_376; // @[Bitwise.scala 71:12]
  wire [9:0] _T_377; // @[Cat.scala 29:58]
  wire [9:0] _T_378; // @[Shift.scala 91:22]
  wire [1:0] _T_379; // @[Shift.scala 92:77]
  wire [7:0] _T_380; // @[Shift.scala 90:30]
  wire [1:0] _T_381; // @[Shift.scala 90:48]
  wire  _T_382; // @[Shift.scala 90:57]
  wire [7:0] _GEN_23; // @[Shift.scala 90:39]
  wire [7:0] _T_383; // @[Shift.scala 90:39]
  wire  _T_384; // @[Shift.scala 12:21]
  wire  _T_385; // @[Shift.scala 12:21]
  wire [1:0] _T_387; // @[Bitwise.scala 71:12]
  wire [9:0] _T_388; // @[Cat.scala 29:58]
  wire [9:0] _T_389; // @[Shift.scala 91:22]
  wire  _T_390; // @[Shift.scala 92:77]
  wire [8:0] _T_391; // @[Shift.scala 90:30]
  wire  _T_392; // @[Shift.scala 90:48]
  wire [8:0] _GEN_24; // @[Shift.scala 90:39]
  wire [8:0] _T_394; // @[Shift.scala 90:39]
  wire  _T_396; // @[Shift.scala 12:21]
  wire [9:0] _T_397; // @[Cat.scala 29:58]
  wire [9:0] _T_398; // @[Shift.scala 91:22]
  wire [9:0] _T_401; // @[Bitwise.scala 71:12]
  wire [9:0] _T_402; // @[Shift.scala 39:10]
  wire  _T_403; // @[convert.scala 55:31]
  wire  _T_404; // @[convert.scala 56:31]
  wire  _T_405; // @[convert.scala 57:31]
  wire  _T_406; // @[convert.scala 58:31]
  wire [6:0] _T_407; // @[convert.scala 59:69]
  wire  _T_408; // @[convert.scala 59:81]
  wire  _T_409; // @[convert.scala 59:50]
  wire  _T_411; // @[convert.scala 60:81]
  wire  _T_412; // @[convert.scala 61:44]
  wire  _T_413; // @[convert.scala 61:52]
  wire  _T_414; // @[convert.scala 61:36]
  wire  _T_415; // @[convert.scala 62:63]
  wire  _T_416; // @[convert.scala 62:103]
  wire  _T_417; // @[convert.scala 62:60]
  wire [6:0] _GEN_25; // @[convert.scala 63:56]
  wire [6:0] _T_420; // @[convert.scala 63:56]
  wire [7:0] _T_421; // @[Cat.scala 29:58]
  wire [7:0] _T_423; // @[Mux.scala 87:16]
  assign _T_1 = io_A[7]; // @[convert.scala 18:24]
  assign _T_2 = io_A[6]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[6:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[5:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[5:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[3:2]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8 != 2'h0; // @[LZD.scala 39:14]
  assign _T_10 = _T_8[1]; // @[LZD.scala 39:21]
  assign _T_11 = _T_8[0]; // @[LZD.scala 39:30]
  assign _T_12 = ~ _T_11; // @[LZD.scala 39:27]
  assign _T_13 = _T_10 | _T_12; // @[LZD.scala 39:25]
  assign _T_14 = {_T_9,_T_13}; // @[Cat.scala 29:58]
  assign _T_15 = _T_7[1:0]; // @[LZD.scala 44:32]
  assign _T_16 = _T_15 != 2'h0; // @[LZD.scala 39:14]
  assign _T_17 = _T_15[1]; // @[LZD.scala 39:21]
  assign _T_18 = _T_15[0]; // @[LZD.scala 39:30]
  assign _T_19 = ~ _T_18; // @[LZD.scala 39:27]
  assign _T_20 = _T_17 | _T_19; // @[LZD.scala 39:25]
  assign _T_21 = {_T_16,_T_20}; // @[Cat.scala 29:58]
  assign _T_22 = _T_14[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22 | _T_23; // @[LZD.scala 49:16]
  assign _T_25 = ~ _T_23; // @[LZD.scala 49:27]
  assign _T_26 = _T_22 | _T_25; // @[LZD.scala 49:25]
  assign _T_27 = _T_14[0:0]; // @[LZD.scala 49:47]
  assign _T_28 = _T_21[0:0]; // @[LZD.scala 49:59]
  assign _T_29 = _T_22 ? _T_27 : _T_28; // @[LZD.scala 49:35]
  assign _T_31 = {_T_24,_T_26,_T_29}; // @[Cat.scala 29:58]
  assign _T_32 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_33 = _T_32 != 2'h0; // @[LZD.scala 39:14]
  assign _T_34 = _T_32[1]; // @[LZD.scala 39:21]
  assign _T_35 = _T_32[0]; // @[LZD.scala 39:30]
  assign _T_36 = ~ _T_35; // @[LZD.scala 39:27]
  assign _T_37 = _T_34 | _T_36; // @[LZD.scala 39:25]
  assign _T_38 = {_T_33,_T_37}; // @[Cat.scala 29:58]
  assign _T_39 = _T_31[2]; // @[Shift.scala 12:21]
  assign _T_41 = _T_31[1:0]; // @[LZD.scala 55:32]
  assign _T_42 = _T_39 ? _T_41 : _T_38; // @[LZD.scala 55:20]
  assign _T_43 = {_T_39,_T_42}; // @[Cat.scala 29:58]
  assign _T_44 = ~ _T_43; // @[convert.scala 21:22]
  assign _T_45 = io_A[4:0]; // @[convert.scala 22:36]
  assign _T_46 = _T_44 < 3'h5; // @[Shift.scala 16:24]
  assign _T_48 = _T_44[2]; // @[Shift.scala 12:21]
  assign _T_49 = _T_45[0:0]; // @[Shift.scala 64:52]
  assign _T_51 = {_T_49,4'h0}; // @[Cat.scala 29:58]
  assign _T_52 = _T_48 ? _T_51 : _T_45; // @[Shift.scala 64:27]
  assign _T_53 = _T_44[1:0]; // @[Shift.scala 66:70]
  assign _T_54 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_55 = _T_52[2:0]; // @[Shift.scala 64:52]
  assign _T_57 = {_T_55,2'h0}; // @[Cat.scala 29:58]
  assign _T_58 = _T_54 ? _T_57 : _T_52; // @[Shift.scala 64:27]
  assign _T_59 = _T_53[0:0]; // @[Shift.scala 66:70]
  assign _T_61 = _T_58[3:0]; // @[Shift.scala 64:52]
  assign _T_62 = {_T_61,1'h0}; // @[Cat.scala 29:58]
  assign _T_63 = _T_59 ? _T_62 : _T_58; // @[Shift.scala 64:27]
  assign _T_64 = _T_46 ? _T_63 : 5'h0; // @[Shift.scala 16:10]
  assign _T_65 = _T_64[4:1]; // @[convert.scala 23:34]
  assign decA_fraction = _T_64[0:0]; // @[convert.scala 24:34]
  assign _T_67 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_69 = _T_3 ? _T_44 : _T_43; // @[convert.scala 25:42]
  assign _T_72 = ~ _T_65; // @[convert.scala 26:67]
  assign _T_73 = _T_1 ? _T_72 : _T_65; // @[convert.scala 26:51]
  assign _T_74 = {_T_67,_T_69,_T_73}; // @[Cat.scala 29:58]
  assign _T_76 = io_A[6:0]; // @[convert.scala 29:56]
  assign _T_77 = _T_76 != 7'h0; // @[convert.scala 29:60]
  assign _T_78 = ~ _T_77; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_78; // @[convert.scala 29:39]
  assign _T_81 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_81 & _T_78; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_74); // @[convert.scala 32:24]
  assign _T_90 = io_B[7]; // @[convert.scala 18:24]
  assign _T_91 = io_B[6]; // @[convert.scala 18:40]
  assign _T_92 = _T_90 ^ _T_91; // @[convert.scala 18:36]
  assign _T_93 = io_B[6:1]; // @[convert.scala 19:24]
  assign _T_94 = io_B[5:0]; // @[convert.scala 19:43]
  assign _T_95 = _T_93 ^ _T_94; // @[convert.scala 19:39]
  assign _T_96 = _T_95[5:2]; // @[LZD.scala 43:32]
  assign _T_97 = _T_96[3:2]; // @[LZD.scala 43:32]
  assign _T_98 = _T_97 != 2'h0; // @[LZD.scala 39:14]
  assign _T_99 = _T_97[1]; // @[LZD.scala 39:21]
  assign _T_100 = _T_97[0]; // @[LZD.scala 39:30]
  assign _T_101 = ~ _T_100; // @[LZD.scala 39:27]
  assign _T_102 = _T_99 | _T_101; // @[LZD.scala 39:25]
  assign _T_103 = {_T_98,_T_102}; // @[Cat.scala 29:58]
  assign _T_104 = _T_96[1:0]; // @[LZD.scala 44:32]
  assign _T_105 = _T_104 != 2'h0; // @[LZD.scala 39:14]
  assign _T_106 = _T_104[1]; // @[LZD.scala 39:21]
  assign _T_107 = _T_104[0]; // @[LZD.scala 39:30]
  assign _T_108 = ~ _T_107; // @[LZD.scala 39:27]
  assign _T_109 = _T_106 | _T_108; // @[LZD.scala 39:25]
  assign _T_110 = {_T_105,_T_109}; // @[Cat.scala 29:58]
  assign _T_111 = _T_103[1]; // @[Shift.scala 12:21]
  assign _T_112 = _T_110[1]; // @[Shift.scala 12:21]
  assign _T_113 = _T_111 | _T_112; // @[LZD.scala 49:16]
  assign _T_114 = ~ _T_112; // @[LZD.scala 49:27]
  assign _T_115 = _T_111 | _T_114; // @[LZD.scala 49:25]
  assign _T_116 = _T_103[0:0]; // @[LZD.scala 49:47]
  assign _T_117 = _T_110[0:0]; // @[LZD.scala 49:59]
  assign _T_118 = _T_111 ? _T_116 : _T_117; // @[LZD.scala 49:35]
  assign _T_120 = {_T_113,_T_115,_T_118}; // @[Cat.scala 29:58]
  assign _T_121 = _T_95[1:0]; // @[LZD.scala 44:32]
  assign _T_122 = _T_121 != 2'h0; // @[LZD.scala 39:14]
  assign _T_123 = _T_121[1]; // @[LZD.scala 39:21]
  assign _T_124 = _T_121[0]; // @[LZD.scala 39:30]
  assign _T_125 = ~ _T_124; // @[LZD.scala 39:27]
  assign _T_126 = _T_123 | _T_125; // @[LZD.scala 39:25]
  assign _T_127 = {_T_122,_T_126}; // @[Cat.scala 29:58]
  assign _T_128 = _T_120[2]; // @[Shift.scala 12:21]
  assign _T_130 = _T_120[1:0]; // @[LZD.scala 55:32]
  assign _T_131 = _T_128 ? _T_130 : _T_127; // @[LZD.scala 55:20]
  assign _T_132 = {_T_128,_T_131}; // @[Cat.scala 29:58]
  assign _T_133 = ~ _T_132; // @[convert.scala 21:22]
  assign _T_134 = io_B[4:0]; // @[convert.scala 22:36]
  assign _T_135 = _T_133 < 3'h5; // @[Shift.scala 16:24]
  assign _T_137 = _T_133[2]; // @[Shift.scala 12:21]
  assign _T_138 = _T_134[0:0]; // @[Shift.scala 64:52]
  assign _T_140 = {_T_138,4'h0}; // @[Cat.scala 29:58]
  assign _T_141 = _T_137 ? _T_140 : _T_134; // @[Shift.scala 64:27]
  assign _T_142 = _T_133[1:0]; // @[Shift.scala 66:70]
  assign _T_143 = _T_142[1]; // @[Shift.scala 12:21]
  assign _T_144 = _T_141[2:0]; // @[Shift.scala 64:52]
  assign _T_146 = {_T_144,2'h0}; // @[Cat.scala 29:58]
  assign _T_147 = _T_143 ? _T_146 : _T_141; // @[Shift.scala 64:27]
  assign _T_148 = _T_142[0:0]; // @[Shift.scala 66:70]
  assign _T_150 = _T_147[3:0]; // @[Shift.scala 64:52]
  assign _T_151 = {_T_150,1'h0}; // @[Cat.scala 29:58]
  assign _T_152 = _T_148 ? _T_151 : _T_147; // @[Shift.scala 64:27]
  assign _T_153 = _T_135 ? _T_152 : 5'h0; // @[Shift.scala 16:10]
  assign _T_154 = _T_153[4:1]; // @[convert.scala 23:34]
  assign decB_fraction = _T_153[0:0]; // @[convert.scala 24:34]
  assign _T_156 = _T_92 == 1'h0; // @[convert.scala 25:26]
  assign _T_158 = _T_92 ? _T_133 : _T_132; // @[convert.scala 25:42]
  assign _T_161 = ~ _T_154; // @[convert.scala 26:67]
  assign _T_162 = _T_90 ? _T_161 : _T_154; // @[convert.scala 26:51]
  assign _T_163 = {_T_156,_T_158,_T_162}; // @[Cat.scala 29:58]
  assign _T_165 = io_B[6:0]; // @[convert.scala 29:56]
  assign _T_166 = _T_165 != 7'h0; // @[convert.scala 29:60]
  assign _T_167 = ~ _T_166; // @[convert.scala 29:41]
  assign decB_isNaR = _T_90 & _T_167; // @[convert.scala 29:39]
  assign _T_170 = _T_90 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_170 & _T_167; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_163); // @[convert.scala 32:24]
  assign _T_179 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_180 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_179,_T_180,decA_fraction,3'h0}; // @[Cat.scala 29:58]
  assign _T_183 = ~ _T_90; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_90,_T_183,decB_fraction,5'h0}; // @[Cat.scala 29:58]
  assign _T_186 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_186 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_187 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_188 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_189 = _T_188 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_190 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_191 = decA_isZero & _T_190; // @[PositDivisionSqrt.scala 94:43]
  assign _T_192 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_193 = _T_191 & _T_192; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_194 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_195 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_194 & _T_195; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_194 & _T_81; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_198 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_198; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 3'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 3'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_199 = sigX_Z[7]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_200 = sigX_Z[5]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_199 ^ _T_200; // @[PositDivisionSqrt.scala 113:50]
  assign _T_201 = cycleNum == 3'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_201 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_202 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_203 = _T_202 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_204 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_205 = entering & _T_204; // @[PositDivisionSqrt.scala 117:30]
  assign _T_207 = io_sqrtOp ? 4'h6 : 4'h8; // @[PositDivisionSqrt.scala 119:26]
  assign _T_208 = entering_normalCase ? _T_207 : 4'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{3'd0}, _T_205}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_209 = _GEN_9 | _T_208; // @[PositDivisionSqrt.scala 117:64]
  assign _T_211 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_212 = _T_202 & _T_211; // @[PositDivisionSqrt.scala 123:27]
  assign _T_214 = cycleNum - 3'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_215 = _T_212 ? _T_214 : 3'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _GEN_10 = {{1'd0}, _T_215}; // @[PositDivisionSqrt.scala 122:64]
  assign _T_216 = _T_209 | _GEN_10; // @[PositDivisionSqrt.scala 122:64]
  assign _T_218 = _T_202 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_11 = {{3'd0}, _T_218}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_220 = _T_216 | _GEN_11; // @[PositDivisionSqrt.scala 123:64]
  assign _GEN_0 = _T_203 ? _T_220 : {{1'd0}, cycleNum}; // @[PositDivisionSqrt.scala 116:29]
  assign _T_221 = decA_scale[7:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_223 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_224 = entering_normalCase & _T_223; // @[PositDivisionSqrt.scala 137:28]
  assign _T_225 = 8'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign _T_226 = _T_225[7:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_227 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_228 = ready & _T_227; // @[PositDivisionSqrt.scala 148:23]
  assign _T_229 = _T_228 ? sigA_S : 8'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_230 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_231 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_232 = _T_231[7:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_233 = _T_230 ? _T_232 : 8'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_234 = _T_229 | _T_233; // @[PositDivisionSqrt.scala 148:66]
  assign _T_235 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_236 = _T_235 ? rem_Z : 8'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_234 | _T_236; // @[PositDivisionSqrt.scala 149:66]
  assign _T_238 = ready & _T_223; // @[PositDivisionSqrt.scala 152:29]
  assign _T_239 = _T_238 ? sigB_S : 8'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_240 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_241 = _T_240 ? 5'h10 : 5'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_12 = {{3'd0}, _T_241}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_242 = _T_239 | _GEN_12; // @[PositDivisionSqrt.scala 152:93]
  assign _T_244 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_245 = _T_235 & _T_244; // @[PositDivisionSqrt.scala 154:30]
  assign _T_246 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_249 = {signB_Z,_T_246,fractB_Z,5'h0}; // @[Cat.scala 29:58]
  assign _T_250 = _T_245 ? _T_249 : 8'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_251 = _T_242 | _T_250; // @[PositDivisionSqrt.scala 153:93]
  assign _T_253 = _T_235 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_254 = rem[7:7]; // @[PositDivisionSqrt.scala 156:83]
  assign _T_256 = _T_254 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign bitMask = {{1'd0}, _T_226}; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  assign _GEN_13 = {{3'd0}, _T_256}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_257 = bitMask & _GEN_13; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_14 = {{1'd0}, _T_257}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_258 = sigX_Z | _GEN_14; // @[PositDivisionSqrt.scala 155:51]
  assign _T_259 = bitMask[6:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_15 = {{2'd0}, _T_259}; // @[PositDivisionSqrt.scala 156:89]
  assign _T_260 = _T_258 | _GEN_15; // @[PositDivisionSqrt.scala 156:89]
  assign _T_261 = _T_253 ? _T_260 : 8'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_251 | _T_261; // @[PositDivisionSqrt.scala 154:93]
  assign _T_263 = trialTerm[7:7]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_264 = _T_254 ^ _T_263; // @[PositDivisionSqrt.scala 162:40]
  assign _T_267 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_269 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_270 = _T_264 ? _T_267 : _T_269; // @[PositDivisionSqrt.scala 161:92]
  assign _T_275 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_276 = _T_275[7:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_278 = _T_276 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_282 = _T_276 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_283 = _T_264 ? _T_278 : _T_282; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_270 : _T_283; // @[PositDivisionSqrt.scala 159:27]
  assign _T_284 = trialRem != 8'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_284 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_285 = rem != 8'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_285 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_287 = trialRem[7:7]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_288 = _T_263 ^ _T_287; // @[PositDivisionSqrt.scala 176:49]
  assign _T_289 = ~ _T_288; // @[PositDivisionSqrt.scala 176:29]
  assign _T_290 = sigX_Z[7:7]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_291 = ~ _T_290; // @[PositDivisionSqrt.scala 178:49]
  assign _T_293 = remIsZero ? _T_290 : _T_289; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_291 : _T_293; // @[Mux.scala 87:16]
  assign _T_294 = cycleNum > 3'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_295 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_296 = _T_294 & _T_295; // @[PositDivisionSqrt.scala 183:48]
  assign _T_297 = entering_normalCase | _T_296; // @[PositDivisionSqrt.scala 183:28]
  assign _T_300 = _T_235 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_301 = entering_normalCase | _T_300; // @[PositDivisionSqrt.scala 187:28]
  assign _T_304 = {newBit, 7'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_305 = _T_238 ? _T_304 : 8'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_307 = _T_240 ? 6'h20 : 6'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_16 = {{2'd0}, _T_307}; // @[PositDivisionSqrt.scala 188:78]
  assign _T_308 = _T_305 | _GEN_16; // @[PositDivisionSqrt.scala 188:78]
  assign _GEN_17 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_310 = sigX_Z | _GEN_17; // @[PositDivisionSqrt.scala 190:47]
  assign _T_311 = _T_235 ? _T_310 : 8'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_312 = _T_308 | _T_311; // @[PositDivisionSqrt.scala 189:78]
  assign _T_314 = {_T_290, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_314 : {{1'd0}, _T_290}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_18 = {{6'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_18; // @[PositDivisionSqrt.scala 197:25]
  assign _T_317 = realSigX[4]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_318 = realSigX[3]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_317 : _T_318; // @[PositDivisionSqrt.scala 198:21]
  assign _T_319 = realSigX[7]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_320 = realSigX[5]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_321 = _T_319 ^ _T_320; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_321; // @[PositDivisionSqrt.scala 205:23]
  assign notNeedSubTwo = _T_319 ^ _T_317; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_324 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_324; // @[PositDivisionSqrt.scala 208:36]
  assign _T_325 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_326 = {1'b0,$signed(_T_325)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_19 = {{6{_T_326[2]}},_T_326}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_328 = $signed(scale_Z) - $signed(_GEN_19); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_328); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-9'sh61); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(9'sh60); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[7:7]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_330 = underflow ? $signed(-9'sh61) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_331 = overflow ? $signed(9'sh60) : $signed(_T_330); // @[Mux.scala 87:16]
  assign _T_332 = realSigX[3:1]; // @[PositDivisionSqrt.scala 224:48]
  assign _T_333 = realSigX[2:0]; // @[PositDivisionSqrt.scala 224:64]
  assign decQ_grs = scaleNotChange ? _T_332 : _T_333; // @[PositDivisionSqrt.scala 224:23]
  assign outValid = cycleNum == 3'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_20 = _T_331[7:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_20); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_339 = decQ_scale[3:0]; // @[convert.scala 46:61]
  assign _T_340 = ~ _T_339; // @[convert.scala 46:52]
  assign _T_342 = decQ_sign ? _T_340 : _T_339; // @[convert.scala 46:42]
  assign _T_343 = decQ_scale[7:4]; // @[convert.scala 48:34]
  assign _T_344 = _T_343[3:3]; // @[convert.scala 49:36]
  assign _T_346 = ~ _T_343; // @[convert.scala 50:36]
  assign _T_347 = $signed(_T_346); // @[convert.scala 50:36]
  assign _T_348 = _T_344 ? $signed(_T_347) : $signed(_T_343); // @[convert.scala 50:28]
  assign _T_349 = _T_344 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_350 = ~ _T_349; // @[convert.scala 52:43]
  assign _T_354 = {_T_350,_T_349,_T_342,realFrac,decQ_grs}; // @[Cat.scala 29:58]
  assign _T_355 = $unsigned(_T_348); // @[Shift.scala 39:17]
  assign _T_356 = _T_355 < 4'ha; // @[Shift.scala 39:24]
  assign _T_358 = _T_354[9:8]; // @[Shift.scala 90:30]
  assign _T_359 = _T_354[7:0]; // @[Shift.scala 90:48]
  assign _T_360 = _T_359 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{1'd0}, _T_360}; // @[Shift.scala 90:39]
  assign _T_361 = _T_358 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_362 = _T_355[3]; // @[Shift.scala 12:21]
  assign _T_363 = _T_354[9]; // @[Shift.scala 12:21]
  assign _T_365 = _T_363 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_366 = {_T_365,_T_361}; // @[Cat.scala 29:58]
  assign _T_367 = _T_362 ? _T_366 : _T_354; // @[Shift.scala 91:22]
  assign _T_368 = _T_355[2:0]; // @[Shift.scala 92:77]
  assign _T_369 = _T_367[9:4]; // @[Shift.scala 90:30]
  assign _T_370 = _T_367[3:0]; // @[Shift.scala 90:48]
  assign _T_371 = _T_370 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{5'd0}, _T_371}; // @[Shift.scala 90:39]
  assign _T_372 = _T_369 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_373 = _T_368[2]; // @[Shift.scala 12:21]
  assign _T_374 = _T_367[9]; // @[Shift.scala 12:21]
  assign _T_376 = _T_374 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_377 = {_T_376,_T_372}; // @[Cat.scala 29:58]
  assign _T_378 = _T_373 ? _T_377 : _T_367; // @[Shift.scala 91:22]
  assign _T_379 = _T_368[1:0]; // @[Shift.scala 92:77]
  assign _T_380 = _T_378[9:2]; // @[Shift.scala 90:30]
  assign _T_381 = _T_378[1:0]; // @[Shift.scala 90:48]
  assign _T_382 = _T_381 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{7'd0}, _T_382}; // @[Shift.scala 90:39]
  assign _T_383 = _T_380 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_384 = _T_379[1]; // @[Shift.scala 12:21]
  assign _T_385 = _T_378[9]; // @[Shift.scala 12:21]
  assign _T_387 = _T_385 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_388 = {_T_387,_T_383}; // @[Cat.scala 29:58]
  assign _T_389 = _T_384 ? _T_388 : _T_378; // @[Shift.scala 91:22]
  assign _T_390 = _T_379[0:0]; // @[Shift.scala 92:77]
  assign _T_391 = _T_389[9:1]; // @[Shift.scala 90:30]
  assign _T_392 = _T_389[0:0]; // @[Shift.scala 90:48]
  assign _GEN_24 = {{8'd0}, _T_392}; // @[Shift.scala 90:39]
  assign _T_394 = _T_391 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_396 = _T_389[9]; // @[Shift.scala 12:21]
  assign _T_397 = {_T_396,_T_394}; // @[Cat.scala 29:58]
  assign _T_398 = _T_390 ? _T_397 : _T_389; // @[Shift.scala 91:22]
  assign _T_401 = _T_363 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_402 = _T_356 ? _T_398 : _T_401; // @[Shift.scala 39:10]
  assign _T_403 = _T_402[3]; // @[convert.scala 55:31]
  assign _T_404 = _T_402[2]; // @[convert.scala 56:31]
  assign _T_405 = _T_402[1]; // @[convert.scala 57:31]
  assign _T_406 = _T_402[0]; // @[convert.scala 58:31]
  assign _T_407 = _T_402[9:3]; // @[convert.scala 59:69]
  assign _T_408 = _T_407 != 7'h0; // @[convert.scala 59:81]
  assign _T_409 = ~ _T_408; // @[convert.scala 59:50]
  assign _T_411 = _T_407 == 7'h7f; // @[convert.scala 60:81]
  assign _T_412 = _T_403 | _T_405; // @[convert.scala 61:44]
  assign _T_413 = _T_412 | _T_406; // @[convert.scala 61:52]
  assign _T_414 = _T_404 & _T_413; // @[convert.scala 61:36]
  assign _T_415 = ~ _T_411; // @[convert.scala 62:63]
  assign _T_416 = _T_415 & _T_414; // @[convert.scala 62:103]
  assign _T_417 = _T_409 | _T_416; // @[convert.scala 62:60]
  assign _GEN_25 = {{6'd0}, _T_417}; // @[convert.scala 63:56]
  assign _T_420 = _T_407 + _GEN_25; // @[convert.scala 63:56]
  assign _T_421 = {decQ_sign,_T_420}; // @[Cat.scala 29:58]
  assign _T_423 = isZero_Z ? 8'h0 : _T_421; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 3'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_244; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 8'h80 : _T_423; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 3'h0;
    end else begin
      cycleNum <= _GEN_0[2:0];
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_187;
      end else begin
        isNaR_Z <= _T_189;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_193;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_221[6]}},_T_221};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_224) begin
      signB_Z <= _T_90;
    end
    if (_T_224) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_297) begin
      if (ready) begin
        if (_T_264) begin
          rem_Z <= _T_267;
        end else begin
          rem_Z <= _T_269;
        end
      end else begin
        if (_T_264) begin
          rem_Z <= _T_278;
        end else begin
          rem_Z <= _T_282;
        end
      end
    end
    if (_T_301) begin
      sigX_Z <= _T_312;
    end
  end
endmodule
