module PositMulEnc6_0(
  input        clock,
  input        reset,
  input  [9:0] io_sigP,
  input  [3:0] io_decAscale,
  input  [3:0] io_decBscale,
  input        io_decAisNar,
  input        io_decBisNar,
  input        io_decAisZero,
  input        io_decBisZero,
  output [5:0] io_M
);
  wire [1:0] head2; // @[PositMulEnc.scala 24:33]
  wire  _T; // @[PositMulEnc.scala 25:31]
  wire  _T_1; // @[PositMulEnc.scala 25:25]
  wire  _T_2; // @[PositMulEnc.scala 25:42]
  wire  addTwo; // @[PositMulEnc.scala 25:35]
  wire  _T_3; // @[PositMulEnc.scala 27:26]
  wire  _T_4; // @[PositMulEnc.scala 27:55]
  wire  addOne; // @[PositMulEnc.scala 27:46]
  wire [1:0] _T_5; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositMulEnc.scala 28:39]
  wire [6:0] _T_6; // @[PositMulEnc.scala 31:84]
  wire [5:0] _T_7; // @[PositMulEnc.scala 32:84]
  wire [6:0] _T_8; // @[PositMulEnc.scala 32:107]
  wire [6:0] frac; // @[PositMulEnc.scala 29:22]
  wire [4:0] _T_9; // @[PositMulEnc.scala 35:32]
  wire [4:0] _GEN_0; // @[PositMulEnc.scala 35:48]
  wire [4:0] _T_11; // @[PositMulEnc.scala 35:48]
  wire [4:0] mulScale; // @[PositMulEnc.scala 35:48]
  wire  underflow; // @[PositMulEnc.scala 36:28]
  wire  overflow; // @[PositMulEnc.scala 37:28]
  wire  decM_sign; // @[PositMulEnc.scala 40:32]
  wire [4:0] _T_14; // @[Mux.scala 87:16]
  wire [4:0] _T_15; // @[Mux.scala 87:16]
  wire [2:0] decM_fraction; // @[PositMulEnc.scala 48:29]
  wire  decM_isNaR; // @[PositMulEnc.scala 49:33]
  wire  decM_isZero; // @[PositMulEnc.scala 50:34]
  wire [3:0] grsTmp; // @[PositMulEnc.scala 53:30]
  wire [1:0] _T_19; // @[PositMulEnc.scala 56:32]
  wire [1:0] _T_20; // @[PositMulEnc.scala 56:48]
  wire  _T_21; // @[PositMulEnc.scala 56:52]
  wire [3:0] _GEN_1; // @[PositMulEnc.scala 39:23 PositMulEnc.scala 41:17]
  wire [3:0] decM_scale; // @[PositMulEnc.scala 39:23 PositMulEnc.scala 41:17]
  wire  _T_25; // @[convert.scala 49:36]
  wire [3:0] _T_27; // @[convert.scala 50:36]
  wire [3:0] _T_28; // @[convert.scala 50:36]
  wire [3:0] _T_29; // @[convert.scala 50:28]
  wire  _T_30; // @[convert.scala 51:31]
  wire  _T_31; // @[convert.scala 53:34]
  wire [7:0] _T_34; // @[Cat.scala 29:58]
  wire [3:0] _T_35; // @[Shift.scala 39:17]
  wire  _T_36; // @[Shift.scala 39:24]
  wire [2:0] _T_37; // @[Shift.scala 40:44]
  wire [3:0] _T_38; // @[Shift.scala 90:30]
  wire [3:0] _T_39; // @[Shift.scala 90:48]
  wire  _T_40; // @[Shift.scala 90:57]
  wire [3:0] _GEN_2; // @[Shift.scala 90:39]
  wire [3:0] _T_41; // @[Shift.scala 90:39]
  wire  _T_42; // @[Shift.scala 12:21]
  wire  _T_43; // @[Shift.scala 12:21]
  wire [3:0] _T_45; // @[Bitwise.scala 71:12]
  wire [7:0] _T_46; // @[Cat.scala 29:58]
  wire [7:0] _T_47; // @[Shift.scala 91:22]
  wire [1:0] _T_48; // @[Shift.scala 92:77]
  wire [5:0] _T_49; // @[Shift.scala 90:30]
  wire [1:0] _T_50; // @[Shift.scala 90:48]
  wire  _T_51; // @[Shift.scala 90:57]
  wire [5:0] _GEN_3; // @[Shift.scala 90:39]
  wire [5:0] _T_52; // @[Shift.scala 90:39]
  wire  _T_53; // @[Shift.scala 12:21]
  wire  _T_54; // @[Shift.scala 12:21]
  wire [1:0] _T_56; // @[Bitwise.scala 71:12]
  wire [7:0] _T_57; // @[Cat.scala 29:58]
  wire [7:0] _T_58; // @[Shift.scala 91:22]
  wire  _T_59; // @[Shift.scala 92:77]
  wire [6:0] _T_60; // @[Shift.scala 90:30]
  wire  _T_61; // @[Shift.scala 90:48]
  wire [6:0] _GEN_4; // @[Shift.scala 90:39]
  wire [6:0] _T_63; // @[Shift.scala 90:39]
  wire  _T_65; // @[Shift.scala 12:21]
  wire [7:0] _T_66; // @[Cat.scala 29:58]
  wire [7:0] _T_67; // @[Shift.scala 91:22]
  wire [7:0] _T_70; // @[Bitwise.scala 71:12]
  wire [7:0] _T_71; // @[Shift.scala 39:10]
  wire  _T_72; // @[convert.scala 55:31]
  wire  _T_73; // @[convert.scala 56:31]
  wire  _T_74; // @[convert.scala 57:31]
  wire  _T_75; // @[convert.scala 58:31]
  wire [4:0] _T_76; // @[convert.scala 59:69]
  wire  _T_77; // @[convert.scala 59:81]
  wire  _T_78; // @[convert.scala 59:50]
  wire  _T_80; // @[convert.scala 60:81]
  wire  _T_81; // @[convert.scala 61:44]
  wire  _T_82; // @[convert.scala 61:52]
  wire  _T_83; // @[convert.scala 61:36]
  wire  _T_84; // @[convert.scala 62:63]
  wire  _T_85; // @[convert.scala 62:103]
  wire  _T_86; // @[convert.scala 62:60]
  wire [4:0] _GEN_5; // @[convert.scala 63:56]
  wire [4:0] _T_89; // @[convert.scala 63:56]
  wire [5:0] _T_90; // @[Cat.scala 29:58]
  wire [5:0] _T_92; // @[Mux.scala 87:16]
  assign head2 = io_sigP[9:8]; // @[PositMulEnc.scala 24:33]
  assign _T = head2[1]; // @[PositMulEnc.scala 25:31]
  assign _T_1 = ~ _T; // @[PositMulEnc.scala 25:25]
  assign _T_2 = head2[0]; // @[PositMulEnc.scala 25:42]
  assign addTwo = _T_1 & _T_2; // @[PositMulEnc.scala 25:35]
  assign _T_3 = io_sigP[9]; // @[PositMulEnc.scala 27:26]
  assign _T_4 = io_sigP[7]; // @[PositMulEnc.scala 27:55]
  assign addOne = _T_3 ^ _T_4; // @[PositMulEnc.scala 27:46]
  assign _T_5 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_5)}; // @[PositMulEnc.scala 28:39]
  assign _T_6 = io_sigP[6:0]; // @[PositMulEnc.scala 31:84]
  assign _T_7 = io_sigP[5:0]; // @[PositMulEnc.scala 32:84]
  assign _T_8 = {_T_7, 1'h0}; // @[PositMulEnc.scala 32:107]
  assign frac = addOne ? _T_6 : _T_8; // @[PositMulEnc.scala 29:22]
  assign _T_9 = $signed(io_decAscale) + $signed(io_decBscale); // @[PositMulEnc.scala 35:32]
  assign _GEN_0 = {{2{expBias[2]}},expBias}; // @[PositMulEnc.scala 35:48]
  assign _T_11 = $signed(_T_9) + $signed(_GEN_0); // @[PositMulEnc.scala 35:48]
  assign mulScale = $signed(_T_11); // @[PositMulEnc.scala 35:48]
  assign underflow = $signed(mulScale) < $signed(-5'sh5); // @[PositMulEnc.scala 36:28]
  assign overflow = $signed(mulScale) > $signed(5'sh4); // @[PositMulEnc.scala 37:28]
  assign decM_sign = io_sigP[9:9]; // @[PositMulEnc.scala 40:32]
  assign _T_14 = underflow ? $signed(-5'sh5) : $signed(mulScale); // @[Mux.scala 87:16]
  assign _T_15 = overflow ? $signed(5'sh4) : $signed(_T_14); // @[Mux.scala 87:16]
  assign decM_fraction = frac[6:4]; // @[PositMulEnc.scala 48:29]
  assign decM_isNaR = io_decAisNar | io_decBisNar; // @[PositMulEnc.scala 49:33]
  assign decM_isZero = io_decAisZero | io_decBisZero; // @[PositMulEnc.scala 50:34]
  assign grsTmp = frac[3:0]; // @[PositMulEnc.scala 53:30]
  assign _T_19 = grsTmp[3:2]; // @[PositMulEnc.scala 56:32]
  assign _T_20 = grsTmp[1:0]; // @[PositMulEnc.scala 56:48]
  assign _T_21 = _T_20 != 2'h0; // @[PositMulEnc.scala 56:52]
  assign _GEN_1 = _T_15[3:0]; // @[PositMulEnc.scala 39:23 PositMulEnc.scala 41:17]
  assign decM_scale = $signed(_GEN_1); // @[PositMulEnc.scala 39:23 PositMulEnc.scala 41:17]
  assign _T_25 = decM_scale[3:3]; // @[convert.scala 49:36]
  assign _T_27 = ~ decM_scale; // @[convert.scala 50:36]
  assign _T_28 = $signed(_T_27); // @[convert.scala 50:36]
  assign _T_29 = _T_25 ? $signed(_T_28) : $signed(decM_scale); // @[convert.scala 50:28]
  assign _T_30 = _T_25 ^ decM_sign; // @[convert.scala 51:31]
  assign _T_31 = ~ _T_30; // @[convert.scala 53:34]
  assign _T_34 = {_T_31,_T_30,decM_fraction,_T_19,_T_21}; // @[Cat.scala 29:58]
  assign _T_35 = $unsigned(_T_29); // @[Shift.scala 39:17]
  assign _T_36 = _T_35 < 4'h8; // @[Shift.scala 39:24]
  assign _T_37 = _T_29[2:0]; // @[Shift.scala 40:44]
  assign _T_38 = _T_34[7:4]; // @[Shift.scala 90:30]
  assign _T_39 = _T_34[3:0]; // @[Shift.scala 90:48]
  assign _T_40 = _T_39 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{3'd0}, _T_40}; // @[Shift.scala 90:39]
  assign _T_41 = _T_38 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_42 = _T_37[2]; // @[Shift.scala 12:21]
  assign _T_43 = _T_34[7]; // @[Shift.scala 12:21]
  assign _T_45 = _T_43 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_46 = {_T_45,_T_41}; // @[Cat.scala 29:58]
  assign _T_47 = _T_42 ? _T_46 : _T_34; // @[Shift.scala 91:22]
  assign _T_48 = _T_37[1:0]; // @[Shift.scala 92:77]
  assign _T_49 = _T_47[7:2]; // @[Shift.scala 90:30]
  assign _T_50 = _T_47[1:0]; // @[Shift.scala 90:48]
  assign _T_51 = _T_50 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_3 = {{5'd0}, _T_51}; // @[Shift.scala 90:39]
  assign _T_52 = _T_49 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_53 = _T_48[1]; // @[Shift.scala 12:21]
  assign _T_54 = _T_47[7]; // @[Shift.scala 12:21]
  assign _T_56 = _T_54 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_57 = {_T_56,_T_52}; // @[Cat.scala 29:58]
  assign _T_58 = _T_53 ? _T_57 : _T_47; // @[Shift.scala 91:22]
  assign _T_59 = _T_48[0:0]; // @[Shift.scala 92:77]
  assign _T_60 = _T_58[7:1]; // @[Shift.scala 90:30]
  assign _T_61 = _T_58[0:0]; // @[Shift.scala 90:48]
  assign _GEN_4 = {{6'd0}, _T_61}; // @[Shift.scala 90:39]
  assign _T_63 = _T_60 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_65 = _T_58[7]; // @[Shift.scala 12:21]
  assign _T_66 = {_T_65,_T_63}; // @[Cat.scala 29:58]
  assign _T_67 = _T_59 ? _T_66 : _T_58; // @[Shift.scala 91:22]
  assign _T_70 = _T_43 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_71 = _T_36 ? _T_67 : _T_70; // @[Shift.scala 39:10]
  assign _T_72 = _T_71[3]; // @[convert.scala 55:31]
  assign _T_73 = _T_71[2]; // @[convert.scala 56:31]
  assign _T_74 = _T_71[1]; // @[convert.scala 57:31]
  assign _T_75 = _T_71[0]; // @[convert.scala 58:31]
  assign _T_76 = _T_71[7:3]; // @[convert.scala 59:69]
  assign _T_77 = _T_76 != 5'h0; // @[convert.scala 59:81]
  assign _T_78 = ~ _T_77; // @[convert.scala 59:50]
  assign _T_80 = _T_76 == 5'h1f; // @[convert.scala 60:81]
  assign _T_81 = _T_72 | _T_74; // @[convert.scala 61:44]
  assign _T_82 = _T_81 | _T_75; // @[convert.scala 61:52]
  assign _T_83 = _T_73 & _T_82; // @[convert.scala 61:36]
  assign _T_84 = ~ _T_80; // @[convert.scala 62:63]
  assign _T_85 = _T_84 & _T_83; // @[convert.scala 62:103]
  assign _T_86 = _T_78 | _T_85; // @[convert.scala 62:60]
  assign _GEN_5 = {{4'd0}, _T_86}; // @[convert.scala 63:56]
  assign _T_89 = _T_76 + _GEN_5; // @[convert.scala 63:56]
  assign _T_90 = {decM_sign,_T_89}; // @[Cat.scala 29:58]
  assign _T_92 = decM_isZero ? 6'h0 : _T_90; // @[Mux.scala 87:16]
  assign io_M = decM_isNaR ? 6'h20 : _T_92; // @[PositMulEnc.scala 64:8]
endmodule
