module FMA_Dec6_0(
  input        clock,
  input        reset,
  input  [5:0] io_A,
  input  [5:0] io_B,
  input  [5:0] io_C,
  output [4:0] io_sigA,
  output [4:0] io_sigB,
  output       io_outIsNaR,
  output       io_Csign,
  output       io_CisNar,
  output       io_CisZero,
  output [2:0] io_Cfrac,
  output [3:0] io_Ascale,
  output [3:0] io_Bscale,
  output [3:0] io_Cscale
);
  wire [6:0] _T_2; // @[FMA_Dec.scala 38:46]
  wire [5:0] realA; // @[FMA_Dec.scala 38:46]
  wire [6:0] _T_5; // @[FMA_Dec.scala 39:46]
  wire [5:0] realC; // @[FMA_Dec.scala 39:46]
  wire  _T_7; // @[convert.scala 18:24]
  wire  _T_8; // @[convert.scala 18:40]
  wire  _T_9; // @[convert.scala 18:36]
  wire [3:0] _T_10; // @[convert.scala 19:24]
  wire [3:0] _T_11; // @[convert.scala 19:43]
  wire [3:0] _T_12; // @[convert.scala 19:39]
  wire [1:0] _T_13; // @[LZD.scala 43:32]
  wire  _T_14; // @[LZD.scala 39:14]
  wire  _T_15; // @[LZD.scala 39:21]
  wire  _T_16; // @[LZD.scala 39:30]
  wire  _T_17; // @[LZD.scala 39:27]
  wire  _T_18; // @[LZD.scala 39:25]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire [1:0] _T_20; // @[LZD.scala 44:32]
  wire  _T_21; // @[LZD.scala 39:14]
  wire  _T_22; // @[LZD.scala 39:21]
  wire  _T_23; // @[LZD.scala 39:30]
  wire  _T_24; // @[LZD.scala 39:27]
  wire  _T_25; // @[LZD.scala 39:25]
  wire [1:0] _T_26; // @[Cat.scala 29:58]
  wire  _T_27; // @[Shift.scala 12:21]
  wire  _T_28; // @[Shift.scala 12:21]
  wire  _T_29; // @[LZD.scala 49:16]
  wire  _T_30; // @[LZD.scala 49:27]
  wire  _T_31; // @[LZD.scala 49:25]
  wire  _T_32; // @[LZD.scala 49:47]
  wire  _T_33; // @[LZD.scala 49:59]
  wire  _T_34; // @[LZD.scala 49:35]
  wire [2:0] _T_36; // @[Cat.scala 29:58]
  wire [2:0] _T_37; // @[convert.scala 21:22]
  wire [2:0] _T_38; // @[convert.scala 22:36]
  wire  _T_39; // @[Shift.scala 16:24]
  wire [1:0] _T_40; // @[Shift.scala 17:37]
  wire  _T_41; // @[Shift.scala 12:21]
  wire  _T_42; // @[Shift.scala 64:52]
  wire [2:0] _T_44; // @[Cat.scala 29:58]
  wire [2:0] _T_45; // @[Shift.scala 64:27]
  wire  _T_46; // @[Shift.scala 66:70]
  wire [1:0] _T_48; // @[Shift.scala 64:52]
  wire [2:0] _T_49; // @[Cat.scala 29:58]
  wire [2:0] _T_50; // @[Shift.scala 64:27]
  wire [2:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_54; // @[convert.scala 25:26]
  wire [2:0] _T_56; // @[convert.scala 25:42]
  wire [3:0] _T_57; // @[Cat.scala 29:58]
  wire [4:0] _T_59; // @[convert.scala 29:56]
  wire  _T_60; // @[convert.scala 29:60]
  wire  _T_61; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_64; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire  _T_73; // @[convert.scala 18:24]
  wire  _T_74; // @[convert.scala 18:40]
  wire  _T_75; // @[convert.scala 18:36]
  wire [3:0] _T_76; // @[convert.scala 19:24]
  wire [3:0] _T_77; // @[convert.scala 19:43]
  wire [3:0] _T_78; // @[convert.scala 19:39]
  wire [1:0] _T_79; // @[LZD.scala 43:32]
  wire  _T_80; // @[LZD.scala 39:14]
  wire  _T_81; // @[LZD.scala 39:21]
  wire  _T_82; // @[LZD.scala 39:30]
  wire  _T_83; // @[LZD.scala 39:27]
  wire  _T_84; // @[LZD.scala 39:25]
  wire [1:0] _T_85; // @[Cat.scala 29:58]
  wire [1:0] _T_86; // @[LZD.scala 44:32]
  wire  _T_87; // @[LZD.scala 39:14]
  wire  _T_88; // @[LZD.scala 39:21]
  wire  _T_89; // @[LZD.scala 39:30]
  wire  _T_90; // @[LZD.scala 39:27]
  wire  _T_91; // @[LZD.scala 39:25]
  wire [1:0] _T_92; // @[Cat.scala 29:58]
  wire  _T_93; // @[Shift.scala 12:21]
  wire  _T_94; // @[Shift.scala 12:21]
  wire  _T_95; // @[LZD.scala 49:16]
  wire  _T_96; // @[LZD.scala 49:27]
  wire  _T_97; // @[LZD.scala 49:25]
  wire  _T_98; // @[LZD.scala 49:47]
  wire  _T_99; // @[LZD.scala 49:59]
  wire  _T_100; // @[LZD.scala 49:35]
  wire [2:0] _T_102; // @[Cat.scala 29:58]
  wire [2:0] _T_103; // @[convert.scala 21:22]
  wire [2:0] _T_104; // @[convert.scala 22:36]
  wire  _T_105; // @[Shift.scala 16:24]
  wire [1:0] _T_106; // @[Shift.scala 17:37]
  wire  _T_107; // @[Shift.scala 12:21]
  wire  _T_108; // @[Shift.scala 64:52]
  wire [2:0] _T_110; // @[Cat.scala 29:58]
  wire [2:0] _T_111; // @[Shift.scala 64:27]
  wire  _T_112; // @[Shift.scala 66:70]
  wire [1:0] _T_114; // @[Shift.scala 64:52]
  wire [2:0] _T_115; // @[Cat.scala 29:58]
  wire [2:0] _T_116; // @[Shift.scala 64:27]
  wire [2:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_120; // @[convert.scala 25:26]
  wire [2:0] _T_122; // @[convert.scala 25:42]
  wire [3:0] _T_123; // @[Cat.scala 29:58]
  wire [4:0] _T_125; // @[convert.scala 29:56]
  wire  _T_126; // @[convert.scala 29:60]
  wire  _T_127; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_130; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire  _T_139; // @[convert.scala 18:24]
  wire  _T_140; // @[convert.scala 18:40]
  wire  _T_141; // @[convert.scala 18:36]
  wire [3:0] _T_142; // @[convert.scala 19:24]
  wire [3:0] _T_143; // @[convert.scala 19:43]
  wire [3:0] _T_144; // @[convert.scala 19:39]
  wire [1:0] _T_145; // @[LZD.scala 43:32]
  wire  _T_146; // @[LZD.scala 39:14]
  wire  _T_147; // @[LZD.scala 39:21]
  wire  _T_148; // @[LZD.scala 39:30]
  wire  _T_149; // @[LZD.scala 39:27]
  wire  _T_150; // @[LZD.scala 39:25]
  wire [1:0] _T_151; // @[Cat.scala 29:58]
  wire [1:0] _T_152; // @[LZD.scala 44:32]
  wire  _T_153; // @[LZD.scala 39:14]
  wire  _T_154; // @[LZD.scala 39:21]
  wire  _T_155; // @[LZD.scala 39:30]
  wire  _T_156; // @[LZD.scala 39:27]
  wire  _T_157; // @[LZD.scala 39:25]
  wire [1:0] _T_158; // @[Cat.scala 29:58]
  wire  _T_159; // @[Shift.scala 12:21]
  wire  _T_160; // @[Shift.scala 12:21]
  wire  _T_161; // @[LZD.scala 49:16]
  wire  _T_162; // @[LZD.scala 49:27]
  wire  _T_163; // @[LZD.scala 49:25]
  wire  _T_164; // @[LZD.scala 49:47]
  wire  _T_165; // @[LZD.scala 49:59]
  wire  _T_166; // @[LZD.scala 49:35]
  wire [2:0] _T_168; // @[Cat.scala 29:58]
  wire [2:0] _T_169; // @[convert.scala 21:22]
  wire [2:0] _T_170; // @[convert.scala 22:36]
  wire  _T_171; // @[Shift.scala 16:24]
  wire [1:0] _T_172; // @[Shift.scala 17:37]
  wire  _T_173; // @[Shift.scala 12:21]
  wire  _T_174; // @[Shift.scala 64:52]
  wire [2:0] _T_176; // @[Cat.scala 29:58]
  wire [2:0] _T_177; // @[Shift.scala 64:27]
  wire  _T_178; // @[Shift.scala 66:70]
  wire [1:0] _T_180; // @[Shift.scala 64:52]
  wire [2:0] _T_181; // @[Cat.scala 29:58]
  wire [2:0] _T_182; // @[Shift.scala 64:27]
  wire  _T_186; // @[convert.scala 25:26]
  wire [2:0] _T_188; // @[convert.scala 25:42]
  wire [3:0] _T_189; // @[Cat.scala 29:58]
  wire [4:0] _T_191; // @[convert.scala 29:56]
  wire  _T_192; // @[convert.scala 29:60]
  wire  _T_193; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_196; // @[convert.scala 30:19]
  wire  _T_204; // @[FMA_Dec.scala 46:30]
  wire  _T_206; // @[FMA_Dec.scala 49:34]
  wire  _T_207; // @[FMA_Dec.scala 49:47]
  wire  _T_208; // @[FMA_Dec.scala 49:45]
  wire [4:0] _T_210; // @[Cat.scala 29:58]
  wire  _T_212; // @[FMA_Dec.scala 50:34]
  wire  _T_213; // @[FMA_Dec.scala 50:47]
  wire  _T_214; // @[FMA_Dec.scala 50:45]
  wire [4:0] _T_216; // @[Cat.scala 29:58]
  assign _T_2 = {{1'd0}, io_A}; // @[FMA_Dec.scala 38:46]
  assign realA = _T_2[5:0]; // @[FMA_Dec.scala 38:46]
  assign _T_5 = {{1'd0}, io_C}; // @[FMA_Dec.scala 39:46]
  assign realC = _T_5[5:0]; // @[FMA_Dec.scala 39:46]
  assign _T_7 = realA[5]; // @[convert.scala 18:24]
  assign _T_8 = realA[4]; // @[convert.scala 18:40]
  assign _T_9 = _T_7 ^ _T_8; // @[convert.scala 18:36]
  assign _T_10 = realA[4:1]; // @[convert.scala 19:24]
  assign _T_11 = realA[3:0]; // @[convert.scala 19:43]
  assign _T_12 = _T_10 ^ _T_11; // @[convert.scala 19:39]
  assign _T_13 = _T_12[3:2]; // @[LZD.scala 43:32]
  assign _T_14 = _T_13 != 2'h0; // @[LZD.scala 39:14]
  assign _T_15 = _T_13[1]; // @[LZD.scala 39:21]
  assign _T_16 = _T_13[0]; // @[LZD.scala 39:30]
  assign _T_17 = ~ _T_16; // @[LZD.scala 39:27]
  assign _T_18 = _T_15 | _T_17; // @[LZD.scala 39:25]
  assign _T_19 = {_T_14,_T_18}; // @[Cat.scala 29:58]
  assign _T_20 = _T_12[1:0]; // @[LZD.scala 44:32]
  assign _T_21 = _T_20 != 2'h0; // @[LZD.scala 39:14]
  assign _T_22 = _T_20[1]; // @[LZD.scala 39:21]
  assign _T_23 = _T_20[0]; // @[LZD.scala 39:30]
  assign _T_24 = ~ _T_23; // @[LZD.scala 39:27]
  assign _T_25 = _T_22 | _T_24; // @[LZD.scala 39:25]
  assign _T_26 = {_T_21,_T_25}; // @[Cat.scala 29:58]
  assign _T_27 = _T_19[1]; // @[Shift.scala 12:21]
  assign _T_28 = _T_26[1]; // @[Shift.scala 12:21]
  assign _T_29 = _T_27 | _T_28; // @[LZD.scala 49:16]
  assign _T_30 = ~ _T_28; // @[LZD.scala 49:27]
  assign _T_31 = _T_27 | _T_30; // @[LZD.scala 49:25]
  assign _T_32 = _T_19[0:0]; // @[LZD.scala 49:47]
  assign _T_33 = _T_26[0:0]; // @[LZD.scala 49:59]
  assign _T_34 = _T_27 ? _T_32 : _T_33; // @[LZD.scala 49:35]
  assign _T_36 = {_T_29,_T_31,_T_34}; // @[Cat.scala 29:58]
  assign _T_37 = ~ _T_36; // @[convert.scala 21:22]
  assign _T_38 = realA[2:0]; // @[convert.scala 22:36]
  assign _T_39 = _T_37 < 3'h3; // @[Shift.scala 16:24]
  assign _T_40 = _T_37[1:0]; // @[Shift.scala 17:37]
  assign _T_41 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_42 = _T_38[0:0]; // @[Shift.scala 64:52]
  assign _T_44 = {_T_42,2'h0}; // @[Cat.scala 29:58]
  assign _T_45 = _T_41 ? _T_44 : _T_38; // @[Shift.scala 64:27]
  assign _T_46 = _T_40[0:0]; // @[Shift.scala 66:70]
  assign _T_48 = _T_45[1:0]; // @[Shift.scala 64:52]
  assign _T_49 = {_T_48,1'h0}; // @[Cat.scala 29:58]
  assign _T_50 = _T_46 ? _T_49 : _T_45; // @[Shift.scala 64:27]
  assign decA_fraction = _T_39 ? _T_50 : 3'h0; // @[Shift.scala 16:10]
  assign _T_54 = _T_9 == 1'h0; // @[convert.scala 25:26]
  assign _T_56 = _T_9 ? _T_37 : _T_36; // @[convert.scala 25:42]
  assign _T_57 = {_T_54,_T_56}; // @[Cat.scala 29:58]
  assign _T_59 = realA[4:0]; // @[convert.scala 29:56]
  assign _T_60 = _T_59 != 5'h0; // @[convert.scala 29:60]
  assign _T_61 = ~ _T_60; // @[convert.scala 29:41]
  assign decA_isNaR = _T_7 & _T_61; // @[convert.scala 29:39]
  assign _T_64 = _T_7 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_64 & _T_61; // @[convert.scala 30:41]
  assign _T_73 = io_B[5]; // @[convert.scala 18:24]
  assign _T_74 = io_B[4]; // @[convert.scala 18:40]
  assign _T_75 = _T_73 ^ _T_74; // @[convert.scala 18:36]
  assign _T_76 = io_B[4:1]; // @[convert.scala 19:24]
  assign _T_77 = io_B[3:0]; // @[convert.scala 19:43]
  assign _T_78 = _T_76 ^ _T_77; // @[convert.scala 19:39]
  assign _T_79 = _T_78[3:2]; // @[LZD.scala 43:32]
  assign _T_80 = _T_79 != 2'h0; // @[LZD.scala 39:14]
  assign _T_81 = _T_79[1]; // @[LZD.scala 39:21]
  assign _T_82 = _T_79[0]; // @[LZD.scala 39:30]
  assign _T_83 = ~ _T_82; // @[LZD.scala 39:27]
  assign _T_84 = _T_81 | _T_83; // @[LZD.scala 39:25]
  assign _T_85 = {_T_80,_T_84}; // @[Cat.scala 29:58]
  assign _T_86 = _T_78[1:0]; // @[LZD.scala 44:32]
  assign _T_87 = _T_86 != 2'h0; // @[LZD.scala 39:14]
  assign _T_88 = _T_86[1]; // @[LZD.scala 39:21]
  assign _T_89 = _T_86[0]; // @[LZD.scala 39:30]
  assign _T_90 = ~ _T_89; // @[LZD.scala 39:27]
  assign _T_91 = _T_88 | _T_90; // @[LZD.scala 39:25]
  assign _T_92 = {_T_87,_T_91}; // @[Cat.scala 29:58]
  assign _T_93 = _T_85[1]; // @[Shift.scala 12:21]
  assign _T_94 = _T_92[1]; // @[Shift.scala 12:21]
  assign _T_95 = _T_93 | _T_94; // @[LZD.scala 49:16]
  assign _T_96 = ~ _T_94; // @[LZD.scala 49:27]
  assign _T_97 = _T_93 | _T_96; // @[LZD.scala 49:25]
  assign _T_98 = _T_85[0:0]; // @[LZD.scala 49:47]
  assign _T_99 = _T_92[0:0]; // @[LZD.scala 49:59]
  assign _T_100 = _T_93 ? _T_98 : _T_99; // @[LZD.scala 49:35]
  assign _T_102 = {_T_95,_T_97,_T_100}; // @[Cat.scala 29:58]
  assign _T_103 = ~ _T_102; // @[convert.scala 21:22]
  assign _T_104 = io_B[2:0]; // @[convert.scala 22:36]
  assign _T_105 = _T_103 < 3'h3; // @[Shift.scala 16:24]
  assign _T_106 = _T_103[1:0]; // @[Shift.scala 17:37]
  assign _T_107 = _T_106[1]; // @[Shift.scala 12:21]
  assign _T_108 = _T_104[0:0]; // @[Shift.scala 64:52]
  assign _T_110 = {_T_108,2'h0}; // @[Cat.scala 29:58]
  assign _T_111 = _T_107 ? _T_110 : _T_104; // @[Shift.scala 64:27]
  assign _T_112 = _T_106[0:0]; // @[Shift.scala 66:70]
  assign _T_114 = _T_111[1:0]; // @[Shift.scala 64:52]
  assign _T_115 = {_T_114,1'h0}; // @[Cat.scala 29:58]
  assign _T_116 = _T_112 ? _T_115 : _T_111; // @[Shift.scala 64:27]
  assign decB_fraction = _T_105 ? _T_116 : 3'h0; // @[Shift.scala 16:10]
  assign _T_120 = _T_75 == 1'h0; // @[convert.scala 25:26]
  assign _T_122 = _T_75 ? _T_103 : _T_102; // @[convert.scala 25:42]
  assign _T_123 = {_T_120,_T_122}; // @[Cat.scala 29:58]
  assign _T_125 = io_B[4:0]; // @[convert.scala 29:56]
  assign _T_126 = _T_125 != 5'h0; // @[convert.scala 29:60]
  assign _T_127 = ~ _T_126; // @[convert.scala 29:41]
  assign decB_isNaR = _T_73 & _T_127; // @[convert.scala 29:39]
  assign _T_130 = _T_73 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_130 & _T_127; // @[convert.scala 30:41]
  assign _T_139 = realC[5]; // @[convert.scala 18:24]
  assign _T_140 = realC[4]; // @[convert.scala 18:40]
  assign _T_141 = _T_139 ^ _T_140; // @[convert.scala 18:36]
  assign _T_142 = realC[4:1]; // @[convert.scala 19:24]
  assign _T_143 = realC[3:0]; // @[convert.scala 19:43]
  assign _T_144 = _T_142 ^ _T_143; // @[convert.scala 19:39]
  assign _T_145 = _T_144[3:2]; // @[LZD.scala 43:32]
  assign _T_146 = _T_145 != 2'h0; // @[LZD.scala 39:14]
  assign _T_147 = _T_145[1]; // @[LZD.scala 39:21]
  assign _T_148 = _T_145[0]; // @[LZD.scala 39:30]
  assign _T_149 = ~ _T_148; // @[LZD.scala 39:27]
  assign _T_150 = _T_147 | _T_149; // @[LZD.scala 39:25]
  assign _T_151 = {_T_146,_T_150}; // @[Cat.scala 29:58]
  assign _T_152 = _T_144[1:0]; // @[LZD.scala 44:32]
  assign _T_153 = _T_152 != 2'h0; // @[LZD.scala 39:14]
  assign _T_154 = _T_152[1]; // @[LZD.scala 39:21]
  assign _T_155 = _T_152[0]; // @[LZD.scala 39:30]
  assign _T_156 = ~ _T_155; // @[LZD.scala 39:27]
  assign _T_157 = _T_154 | _T_156; // @[LZD.scala 39:25]
  assign _T_158 = {_T_153,_T_157}; // @[Cat.scala 29:58]
  assign _T_159 = _T_151[1]; // @[Shift.scala 12:21]
  assign _T_160 = _T_158[1]; // @[Shift.scala 12:21]
  assign _T_161 = _T_159 | _T_160; // @[LZD.scala 49:16]
  assign _T_162 = ~ _T_160; // @[LZD.scala 49:27]
  assign _T_163 = _T_159 | _T_162; // @[LZD.scala 49:25]
  assign _T_164 = _T_151[0:0]; // @[LZD.scala 49:47]
  assign _T_165 = _T_158[0:0]; // @[LZD.scala 49:59]
  assign _T_166 = _T_159 ? _T_164 : _T_165; // @[LZD.scala 49:35]
  assign _T_168 = {_T_161,_T_163,_T_166}; // @[Cat.scala 29:58]
  assign _T_169 = ~ _T_168; // @[convert.scala 21:22]
  assign _T_170 = realC[2:0]; // @[convert.scala 22:36]
  assign _T_171 = _T_169 < 3'h3; // @[Shift.scala 16:24]
  assign _T_172 = _T_169[1:0]; // @[Shift.scala 17:37]
  assign _T_173 = _T_172[1]; // @[Shift.scala 12:21]
  assign _T_174 = _T_170[0:0]; // @[Shift.scala 64:52]
  assign _T_176 = {_T_174,2'h0}; // @[Cat.scala 29:58]
  assign _T_177 = _T_173 ? _T_176 : _T_170; // @[Shift.scala 64:27]
  assign _T_178 = _T_172[0:0]; // @[Shift.scala 66:70]
  assign _T_180 = _T_177[1:0]; // @[Shift.scala 64:52]
  assign _T_181 = {_T_180,1'h0}; // @[Cat.scala 29:58]
  assign _T_182 = _T_178 ? _T_181 : _T_177; // @[Shift.scala 64:27]
  assign _T_186 = _T_141 == 1'h0; // @[convert.scala 25:26]
  assign _T_188 = _T_141 ? _T_169 : _T_168; // @[convert.scala 25:42]
  assign _T_189 = {_T_186,_T_188}; // @[Cat.scala 29:58]
  assign _T_191 = realC[4:0]; // @[convert.scala 29:56]
  assign _T_192 = _T_191 != 5'h0; // @[convert.scala 29:60]
  assign _T_193 = ~ _T_192; // @[convert.scala 29:41]
  assign decC_isNaR = _T_139 & _T_193; // @[convert.scala 29:39]
  assign _T_196 = _T_139 == 1'h0; // @[convert.scala 30:19]
  assign _T_204 = decA_isNaR | decB_isNaR; // @[FMA_Dec.scala 46:30]
  assign _T_206 = ~ _T_7; // @[FMA_Dec.scala 49:34]
  assign _T_207 = ~ decA_isZero; // @[FMA_Dec.scala 49:47]
  assign _T_208 = _T_206 & _T_207; // @[FMA_Dec.scala 49:45]
  assign _T_210 = {_T_7,_T_208,decA_fraction}; // @[Cat.scala 29:58]
  assign _T_212 = ~ _T_73; // @[FMA_Dec.scala 50:34]
  assign _T_213 = ~ decB_isZero; // @[FMA_Dec.scala 50:47]
  assign _T_214 = _T_212 & _T_213; // @[FMA_Dec.scala 50:45]
  assign _T_216 = {_T_73,_T_214,decB_fraction}; // @[Cat.scala 29:58]
  assign io_sigA = $signed(_T_210); // @[FMA_Dec.scala 49:16]
  assign io_sigB = $signed(_T_216); // @[FMA_Dec.scala 50:16]
  assign io_outIsNaR = _T_204 | decC_isNaR; // @[FMA_Dec.scala 46:16]
  assign io_Csign = realC[5]; // @[FMA_Dec.scala 55:12]
  assign io_CisNar = _T_139 & _T_193; // @[FMA_Dec.scala 51:17]
  assign io_CisZero = _T_196 & _T_193; // @[FMA_Dec.scala 52:17]
  assign io_Cfrac = _T_171 ? _T_182 : 3'h0; // @[FMA_Dec.scala 53:17]
  assign io_Ascale = $signed(_T_57); // @[FMA_Dec.scala 47:13]
  assign io_Bscale = $signed(_T_123); // @[FMA_Dec.scala 48:13]
  assign io_Cscale = $signed(_T_189); // @[FMA_Dec.scala 54:16]
endmodule
