module Post_Adder5_1(
  input        clock,
  input        reset,
  input  [6:0] io_signSumSig,
  input  [3:0] io_greaterExp,
  input        io_sumSign,
  output       io_overflow,
  input        io_AisNar,
  input        io_BisNar,
  input        io_AisZero,
  input        io_BisZero,
  output [4:0] io_S
);
  wire [5:0] _T; // @[Post_Adder.scala 26:34]
  wire [5:0] _T_1; // @[Post_Adder.scala 26:72]
  wire [5:0] sumXor; // @[Post_Adder.scala 26:52]
  wire [3:0] _T_2; // @[LZD.scala 43:32]
  wire [1:0] _T_3; // @[LZD.scala 43:32]
  wire  _T_4; // @[LZD.scala 39:14]
  wire  _T_5; // @[LZD.scala 39:21]
  wire  _T_6; // @[LZD.scala 39:30]
  wire  _T_7; // @[LZD.scala 39:27]
  wire  _T_8; // @[LZD.scala 39:25]
  wire [1:0] _T_9; // @[Cat.scala 29:58]
  wire [1:0] _T_10; // @[LZD.scala 44:32]
  wire  _T_11; // @[LZD.scala 39:14]
  wire  _T_12; // @[LZD.scala 39:21]
  wire  _T_13; // @[LZD.scala 39:30]
  wire  _T_14; // @[LZD.scala 39:27]
  wire  _T_15; // @[LZD.scala 39:25]
  wire [1:0] _T_16; // @[Cat.scala 29:58]
  wire  _T_17; // @[Shift.scala 12:21]
  wire  _T_18; // @[Shift.scala 12:21]
  wire  _T_19; // @[LZD.scala 49:16]
  wire  _T_20; // @[LZD.scala 49:27]
  wire  _T_21; // @[LZD.scala 49:25]
  wire  _T_22; // @[LZD.scala 49:47]
  wire  _T_23; // @[LZD.scala 49:59]
  wire  _T_24; // @[LZD.scala 49:35]
  wire [2:0] _T_26; // @[Cat.scala 29:58]
  wire [1:0] _T_27; // @[LZD.scala 44:32]
  wire  _T_28; // @[LZD.scala 39:14]
  wire  _T_29; // @[LZD.scala 39:21]
  wire  _T_30; // @[LZD.scala 39:30]
  wire  _T_31; // @[LZD.scala 39:27]
  wire  _T_32; // @[LZD.scala 39:25]
  wire [1:0] _T_33; // @[Cat.scala 29:58]
  wire  _T_34; // @[Shift.scala 12:21]
  wire [1:0] _T_36; // @[LZD.scala 55:32]
  wire [1:0] _T_37; // @[LZD.scala 55:20]
  wire [2:0] sumLZD; // @[Cat.scala 29:58]
  wire [3:0] _T_38; // @[Cat.scala 29:58]
  wire [3:0] _T_39; // @[Post_Adder.scala 28:37]
  wire [3:0] _T_41; // @[Post_Adder.scala 28:44]
  wire [3:0] scaleBias; // @[Post_Adder.scala 28:44]
  wire [4:0] sumScale; // @[Post_Adder.scala 29:35]
  wire [2:0] normalShift; // @[Post_Adder.scala 31:22]
  wire [4:0] _T_43; // @[Post_Adder.scala 32:39]
  wire  _T_44; // @[Shift.scala 16:24]
  wire  _T_46; // @[Shift.scala 12:21]
  wire  _T_47; // @[Shift.scala 64:52]
  wire [4:0] _T_49; // @[Cat.scala 29:58]
  wire [4:0] _T_50; // @[Shift.scala 64:27]
  wire [1:0] _T_51; // @[Shift.scala 66:70]
  wire  _T_52; // @[Shift.scala 12:21]
  wire [2:0] _T_53; // @[Shift.scala 64:52]
  wire [4:0] _T_55; // @[Cat.scala 29:58]
  wire [4:0] _T_56; // @[Shift.scala 64:27]
  wire  _T_57; // @[Shift.scala 66:70]
  wire [3:0] _T_59; // @[Shift.scala 64:52]
  wire [4:0] _T_60; // @[Cat.scala 29:58]
  wire [4:0] _T_61; // @[Shift.scala 64:27]
  wire [4:0] shiftSig; // @[Shift.scala 16:10]
  wire [4:0] _T_62; // @[Post_Adder.scala 44:24]
  wire  decS_fraction; // @[Post_Adder.scala 45:34]
  wire  decS_isNaR; // @[Post_Adder.scala 46:31]
  wire  _T_65; // @[Post_Adder.scala 47:36]
  wire  _T_66; // @[Post_Adder.scala 47:21]
  wire  _T_67; // @[Post_Adder.scala 47:54]
  wire  decS_isZero; // @[Post_Adder.scala 47:40]
  wire [1:0] _T_69; // @[Post_Adder.scala 48:33]
  wire  _T_70; // @[Post_Adder.scala 48:49]
  wire  _T_71; // @[Post_Adder.scala 48:63]
  wire  _T_72; // @[Post_Adder.scala 48:53]
  wire [3:0] _GEN_0; // @[Post_Adder.scala 41:24 Post_Adder.scala 44:18]
  wire [3:0] decS_scale; // @[Post_Adder.scala 41:24 Post_Adder.scala 44:18]
  wire  _T_75; // @[convert.scala 46:61]
  wire  _T_76; // @[convert.scala 46:52]
  wire  _T_78; // @[convert.scala 46:42]
  wire [2:0] _T_79; // @[convert.scala 48:34]
  wire  _T_80; // @[convert.scala 49:36]
  wire [2:0] _T_82; // @[convert.scala 50:36]
  wire [2:0] _T_83; // @[convert.scala 50:36]
  wire [2:0] _T_84; // @[convert.scala 50:28]
  wire  _T_85; // @[convert.scala 51:31]
  wire  _T_86; // @[convert.scala 52:43]
  wire [6:0] _T_90; // @[Cat.scala 29:58]
  wire [2:0] _T_91; // @[Shift.scala 39:17]
  wire  _T_92; // @[Shift.scala 39:24]
  wire [2:0] _T_94; // @[Shift.scala 90:30]
  wire [3:0] _T_95; // @[Shift.scala 90:48]
  wire  _T_96; // @[Shift.scala 90:57]
  wire [2:0] _GEN_1; // @[Shift.scala 90:39]
  wire [2:0] _T_97; // @[Shift.scala 90:39]
  wire  _T_98; // @[Shift.scala 12:21]
  wire  _T_99; // @[Shift.scala 12:21]
  wire [3:0] _T_101; // @[Bitwise.scala 71:12]
  wire [6:0] _T_102; // @[Cat.scala 29:58]
  wire [6:0] _T_103; // @[Shift.scala 91:22]
  wire [1:0] _T_104; // @[Shift.scala 92:77]
  wire [4:0] _T_105; // @[Shift.scala 90:30]
  wire [1:0] _T_106; // @[Shift.scala 90:48]
  wire  _T_107; // @[Shift.scala 90:57]
  wire [4:0] _GEN_2; // @[Shift.scala 90:39]
  wire [4:0] _T_108; // @[Shift.scala 90:39]
  wire  _T_109; // @[Shift.scala 12:21]
  wire  _T_110; // @[Shift.scala 12:21]
  wire [1:0] _T_112; // @[Bitwise.scala 71:12]
  wire [6:0] _T_113; // @[Cat.scala 29:58]
  wire [6:0] _T_114; // @[Shift.scala 91:22]
  wire  _T_115; // @[Shift.scala 92:77]
  wire [5:0] _T_116; // @[Shift.scala 90:30]
  wire  _T_117; // @[Shift.scala 90:48]
  wire [5:0] _GEN_3; // @[Shift.scala 90:39]
  wire [5:0] _T_119; // @[Shift.scala 90:39]
  wire  _T_121; // @[Shift.scala 12:21]
  wire [6:0] _T_122; // @[Cat.scala 29:58]
  wire [6:0] _T_123; // @[Shift.scala 91:22]
  wire [6:0] _T_126; // @[Bitwise.scala 71:12]
  wire [6:0] _T_127; // @[Shift.scala 39:10]
  wire  _T_128; // @[convert.scala 55:31]
  wire  _T_129; // @[convert.scala 56:31]
  wire  _T_130; // @[convert.scala 57:31]
  wire  _T_131; // @[convert.scala 58:31]
  wire [3:0] _T_132; // @[convert.scala 59:69]
  wire  _T_133; // @[convert.scala 59:81]
  wire  _T_134; // @[convert.scala 59:50]
  wire  _T_136; // @[convert.scala 60:81]
  wire  _T_137; // @[convert.scala 61:44]
  wire  _T_138; // @[convert.scala 61:52]
  wire  _T_139; // @[convert.scala 61:36]
  wire  _T_140; // @[convert.scala 62:63]
  wire  _T_141; // @[convert.scala 62:103]
  wire  _T_142; // @[convert.scala 62:60]
  wire [3:0] _GEN_4; // @[convert.scala 63:56]
  wire [3:0] _T_145; // @[convert.scala 63:56]
  wire [4:0] _T_146; // @[Cat.scala 29:58]
  wire [4:0] _T_148; // @[Mux.scala 87:16]
  assign _T = io_signSumSig[6:1]; // @[Post_Adder.scala 26:34]
  assign _T_1 = io_signSumSig[5:0]; // @[Post_Adder.scala 26:72]
  assign sumXor = _T ^ _T_1; // @[Post_Adder.scala 26:52]
  assign _T_2 = sumXor[5:2]; // @[LZD.scala 43:32]
  assign _T_3 = _T_2[3:2]; // @[LZD.scala 43:32]
  assign _T_4 = _T_3 != 2'h0; // @[LZD.scala 39:14]
  assign _T_5 = _T_3[1]; // @[LZD.scala 39:21]
  assign _T_6 = _T_3[0]; // @[LZD.scala 39:30]
  assign _T_7 = ~ _T_6; // @[LZD.scala 39:27]
  assign _T_8 = _T_5 | _T_7; // @[LZD.scala 39:25]
  assign _T_9 = {_T_4,_T_8}; // @[Cat.scala 29:58]
  assign _T_10 = _T_2[1:0]; // @[LZD.scala 44:32]
  assign _T_11 = _T_10 != 2'h0; // @[LZD.scala 39:14]
  assign _T_12 = _T_10[1]; // @[LZD.scala 39:21]
  assign _T_13 = _T_10[0]; // @[LZD.scala 39:30]
  assign _T_14 = ~ _T_13; // @[LZD.scala 39:27]
  assign _T_15 = _T_12 | _T_14; // @[LZD.scala 39:25]
  assign _T_16 = {_T_11,_T_15}; // @[Cat.scala 29:58]
  assign _T_17 = _T_9[1]; // @[Shift.scala 12:21]
  assign _T_18 = _T_16[1]; // @[Shift.scala 12:21]
  assign _T_19 = _T_17 | _T_18; // @[LZD.scala 49:16]
  assign _T_20 = ~ _T_18; // @[LZD.scala 49:27]
  assign _T_21 = _T_17 | _T_20; // @[LZD.scala 49:25]
  assign _T_22 = _T_9[0:0]; // @[LZD.scala 49:47]
  assign _T_23 = _T_16[0:0]; // @[LZD.scala 49:59]
  assign _T_24 = _T_17 ? _T_22 : _T_23; // @[LZD.scala 49:35]
  assign _T_26 = {_T_19,_T_21,_T_24}; // @[Cat.scala 29:58]
  assign _T_27 = sumXor[1:0]; // @[LZD.scala 44:32]
  assign _T_28 = _T_27 != 2'h0; // @[LZD.scala 39:14]
  assign _T_29 = _T_27[1]; // @[LZD.scala 39:21]
  assign _T_30 = _T_27[0]; // @[LZD.scala 39:30]
  assign _T_31 = ~ _T_30; // @[LZD.scala 39:27]
  assign _T_32 = _T_29 | _T_31; // @[LZD.scala 39:25]
  assign _T_33 = {_T_28,_T_32}; // @[Cat.scala 29:58]
  assign _T_34 = _T_26[2]; // @[Shift.scala 12:21]
  assign _T_36 = _T_26[1:0]; // @[LZD.scala 55:32]
  assign _T_37 = _T_34 ? _T_36 : _T_33; // @[LZD.scala 55:20]
  assign sumLZD = {_T_34,_T_37}; // @[Cat.scala 29:58]
  assign _T_38 = {1'h1,_T_34,_T_37}; // @[Cat.scala 29:58]
  assign _T_39 = $signed(_T_38); // @[Post_Adder.scala 28:37]
  assign _T_41 = $signed(_T_39) + $signed(4'sh2); // @[Post_Adder.scala 28:44]
  assign scaleBias = $signed(_T_41); // @[Post_Adder.scala 28:44]
  assign sumScale = $signed(io_greaterExp) + $signed(scaleBias); // @[Post_Adder.scala 29:35]
  assign normalShift = ~ sumLZD; // @[Post_Adder.scala 31:22]
  assign _T_43 = io_signSumSig[4:0]; // @[Post_Adder.scala 32:39]
  assign _T_44 = normalShift < 3'h5; // @[Shift.scala 16:24]
  assign _T_46 = normalShift[2]; // @[Shift.scala 12:21]
  assign _T_47 = _T_43[0:0]; // @[Shift.scala 64:52]
  assign _T_49 = {_T_47,4'h0}; // @[Cat.scala 29:58]
  assign _T_50 = _T_46 ? _T_49 : _T_43; // @[Shift.scala 64:27]
  assign _T_51 = normalShift[1:0]; // @[Shift.scala 66:70]
  assign _T_52 = _T_51[1]; // @[Shift.scala 12:21]
  assign _T_53 = _T_50[2:0]; // @[Shift.scala 64:52]
  assign _T_55 = {_T_53,2'h0}; // @[Cat.scala 29:58]
  assign _T_56 = _T_52 ? _T_55 : _T_50; // @[Shift.scala 64:27]
  assign _T_57 = _T_51[0:0]; // @[Shift.scala 66:70]
  assign _T_59 = _T_56[3:0]; // @[Shift.scala 64:52]
  assign _T_60 = {_T_59,1'h0}; // @[Cat.scala 29:58]
  assign _T_61 = _T_57 ? _T_60 : _T_56; // @[Shift.scala 64:27]
  assign shiftSig = _T_44 ? _T_61 : 5'h0; // @[Shift.scala 16:10]
  assign _T_62 = io_overflow ? $signed(5'sh6) : $signed(sumScale); // @[Post_Adder.scala 44:24]
  assign decS_fraction = shiftSig[4:4]; // @[Post_Adder.scala 45:34]
  assign decS_isNaR = io_AisNar | io_BisNar; // @[Post_Adder.scala 46:31]
  assign _T_65 = io_signSumSig != 7'h0; // @[Post_Adder.scala 47:36]
  assign _T_66 = ~ _T_65; // @[Post_Adder.scala 47:21]
  assign _T_67 = io_AisZero & io_BisZero; // @[Post_Adder.scala 47:54]
  assign decS_isZero = _T_66 | _T_67; // @[Post_Adder.scala 47:40]
  assign _T_69 = shiftSig[3:2]; // @[Post_Adder.scala 48:33]
  assign _T_70 = shiftSig[1]; // @[Post_Adder.scala 48:49]
  assign _T_71 = shiftSig[0]; // @[Post_Adder.scala 48:63]
  assign _T_72 = _T_70 | _T_71; // @[Post_Adder.scala 48:53]
  assign _GEN_0 = _T_62[3:0]; // @[Post_Adder.scala 41:24 Post_Adder.scala 44:18]
  assign decS_scale = $signed(_GEN_0); // @[Post_Adder.scala 41:24 Post_Adder.scala 44:18]
  assign _T_75 = decS_scale[0]; // @[convert.scala 46:61]
  assign _T_76 = ~ _T_75; // @[convert.scala 46:52]
  assign _T_78 = io_sumSign ? _T_76 : _T_75; // @[convert.scala 46:42]
  assign _T_79 = decS_scale[3:1]; // @[convert.scala 48:34]
  assign _T_80 = _T_79[2:2]; // @[convert.scala 49:36]
  assign _T_82 = ~ _T_79; // @[convert.scala 50:36]
  assign _T_83 = $signed(_T_82); // @[convert.scala 50:36]
  assign _T_84 = _T_80 ? $signed(_T_83) : $signed(_T_79); // @[convert.scala 50:28]
  assign _T_85 = _T_80 ^ io_sumSign; // @[convert.scala 51:31]
  assign _T_86 = ~ _T_85; // @[convert.scala 52:43]
  assign _T_90 = {_T_86,_T_85,_T_78,decS_fraction,_T_69,_T_72}; // @[Cat.scala 29:58]
  assign _T_91 = $unsigned(_T_84); // @[Shift.scala 39:17]
  assign _T_92 = _T_91 < 3'h7; // @[Shift.scala 39:24]
  assign _T_94 = _T_90[6:4]; // @[Shift.scala 90:30]
  assign _T_95 = _T_90[3:0]; // @[Shift.scala 90:48]
  assign _T_96 = _T_95 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{2'd0}, _T_96}; // @[Shift.scala 90:39]
  assign _T_97 = _T_94 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_98 = _T_91[2]; // @[Shift.scala 12:21]
  assign _T_99 = _T_90[6]; // @[Shift.scala 12:21]
  assign _T_101 = _T_99 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_102 = {_T_101,_T_97}; // @[Cat.scala 29:58]
  assign _T_103 = _T_98 ? _T_102 : _T_90; // @[Shift.scala 91:22]
  assign _T_104 = _T_91[1:0]; // @[Shift.scala 92:77]
  assign _T_105 = _T_103[6:2]; // @[Shift.scala 90:30]
  assign _T_106 = _T_103[1:0]; // @[Shift.scala 90:48]
  assign _T_107 = _T_106 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{4'd0}, _T_107}; // @[Shift.scala 90:39]
  assign _T_108 = _T_105 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_109 = _T_104[1]; // @[Shift.scala 12:21]
  assign _T_110 = _T_103[6]; // @[Shift.scala 12:21]
  assign _T_112 = _T_110 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_113 = {_T_112,_T_108}; // @[Cat.scala 29:58]
  assign _T_114 = _T_109 ? _T_113 : _T_103; // @[Shift.scala 91:22]
  assign _T_115 = _T_104[0:0]; // @[Shift.scala 92:77]
  assign _T_116 = _T_114[6:1]; // @[Shift.scala 90:30]
  assign _T_117 = _T_114[0:0]; // @[Shift.scala 90:48]
  assign _GEN_3 = {{5'd0}, _T_117}; // @[Shift.scala 90:39]
  assign _T_119 = _T_116 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_121 = _T_114[6]; // @[Shift.scala 12:21]
  assign _T_122 = {_T_121,_T_119}; // @[Cat.scala 29:58]
  assign _T_123 = _T_115 ? _T_122 : _T_114; // @[Shift.scala 91:22]
  assign _T_126 = _T_99 ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign _T_127 = _T_92 ? _T_123 : _T_126; // @[Shift.scala 39:10]
  assign _T_128 = _T_127[3]; // @[convert.scala 55:31]
  assign _T_129 = _T_127[2]; // @[convert.scala 56:31]
  assign _T_130 = _T_127[1]; // @[convert.scala 57:31]
  assign _T_131 = _T_127[0]; // @[convert.scala 58:31]
  assign _T_132 = _T_127[6:3]; // @[convert.scala 59:69]
  assign _T_133 = _T_132 != 4'h0; // @[convert.scala 59:81]
  assign _T_134 = ~ _T_133; // @[convert.scala 59:50]
  assign _T_136 = _T_132 == 4'hf; // @[convert.scala 60:81]
  assign _T_137 = _T_128 | _T_130; // @[convert.scala 61:44]
  assign _T_138 = _T_137 | _T_131; // @[convert.scala 61:52]
  assign _T_139 = _T_129 & _T_138; // @[convert.scala 61:36]
  assign _T_140 = ~ _T_136; // @[convert.scala 62:63]
  assign _T_141 = _T_140 & _T_139; // @[convert.scala 62:103]
  assign _T_142 = _T_134 | _T_141; // @[convert.scala 62:60]
  assign _GEN_4 = {{3'd0}, _T_142}; // @[convert.scala 63:56]
  assign _T_145 = _T_132 + _GEN_4; // @[convert.scala 63:56]
  assign _T_146 = {io_sumSign,_T_145}; // @[Cat.scala 29:58]
  assign _T_148 = decS_isZero ? 5'h0 : _T_146; // @[Mux.scala 87:16]
  assign io_overflow = $signed(sumScale) > $signed(5'sh6); // @[Post_Adder.scala 30:18]
  assign io_S = decS_isNaR ? 5'h10 : _T_148; // @[Post_Adder.scala 49:7]
endmodule
