module PositDivSqrter6_2(
  input        clock,
  input        reset,
  output       io_inReady,
  input        io_inValid,
  input        io_sqrtOp,
  input  [5:0] io_A,
  input  [5:0] io_B,
  output       io_diviValid,
  output       io_sqrtValid,
  output       io_invalidExc,
  output [5:0] io_Q
);
  reg [2:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [6:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg  fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [7:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [7:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [3:0] _T_4; // @[convert.scala 19:24]
  wire [3:0] _T_5; // @[convert.scala 19:43]
  wire [3:0] _T_6; // @[convert.scala 19:39]
  wire [1:0] _T_7; // @[LZD.scala 43:32]
  wire  _T_8; // @[LZD.scala 39:14]
  wire  _T_9; // @[LZD.scala 39:21]
  wire  _T_10; // @[LZD.scala 39:30]
  wire  _T_11; // @[LZD.scala 39:27]
  wire  _T_12; // @[LZD.scala 39:25]
  wire [1:0] _T_13; // @[Cat.scala 29:58]
  wire [1:0] _T_14; // @[LZD.scala 44:32]
  wire  _T_15; // @[LZD.scala 39:14]
  wire  _T_16; // @[LZD.scala 39:21]
  wire  _T_17; // @[LZD.scala 39:30]
  wire  _T_18; // @[LZD.scala 39:27]
  wire  _T_19; // @[LZD.scala 39:25]
  wire [1:0] _T_20; // @[Cat.scala 29:58]
  wire  _T_21; // @[Shift.scala 12:21]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[LZD.scala 49:16]
  wire  _T_24; // @[LZD.scala 49:27]
  wire  _T_25; // @[LZD.scala 49:25]
  wire  _T_26; // @[LZD.scala 49:47]
  wire  _T_27; // @[LZD.scala 49:59]
  wire  _T_28; // @[LZD.scala 49:35]
  wire [2:0] _T_30; // @[Cat.scala 29:58]
  wire [2:0] _T_31; // @[convert.scala 21:22]
  wire [2:0] _T_32; // @[convert.scala 22:36]
  wire  _T_33; // @[Shift.scala 16:24]
  wire [1:0] _T_34; // @[Shift.scala 17:37]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[Shift.scala 64:52]
  wire [2:0] _T_38; // @[Cat.scala 29:58]
  wire [2:0] _T_39; // @[Shift.scala 64:27]
  wire  _T_40; // @[Shift.scala 66:70]
  wire [1:0] _T_42; // @[Shift.scala 64:52]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire [2:0] _T_44; // @[Shift.scala 64:27]
  wire [2:0] _T_45; // @[Shift.scala 16:10]
  wire [1:0] _T_46; // @[convert.scala 23:34]
  wire  decA_fraction; // @[convert.scala 24:34]
  wire  _T_48; // @[convert.scala 25:26]
  wire [2:0] _T_50; // @[convert.scala 25:42]
  wire [1:0] _T_53; // @[convert.scala 26:67]
  wire [1:0] _T_54; // @[convert.scala 26:51]
  wire [5:0] _T_55; // @[Cat.scala 29:58]
  wire [4:0] _T_57; // @[convert.scala 29:56]
  wire  _T_58; // @[convert.scala 29:60]
  wire  _T_59; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_62; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_71; // @[convert.scala 18:24]
  wire  _T_72; // @[convert.scala 18:40]
  wire  _T_73; // @[convert.scala 18:36]
  wire [3:0] _T_74; // @[convert.scala 19:24]
  wire [3:0] _T_75; // @[convert.scala 19:43]
  wire [3:0] _T_76; // @[convert.scala 19:39]
  wire [1:0] _T_77; // @[LZD.scala 43:32]
  wire  _T_78; // @[LZD.scala 39:14]
  wire  _T_79; // @[LZD.scala 39:21]
  wire  _T_80; // @[LZD.scala 39:30]
  wire  _T_81; // @[LZD.scala 39:27]
  wire  _T_82; // @[LZD.scala 39:25]
  wire [1:0] _T_83; // @[Cat.scala 29:58]
  wire [1:0] _T_84; // @[LZD.scala 44:32]
  wire  _T_85; // @[LZD.scala 39:14]
  wire  _T_86; // @[LZD.scala 39:21]
  wire  _T_87; // @[LZD.scala 39:30]
  wire  _T_88; // @[LZD.scala 39:27]
  wire  _T_89; // @[LZD.scala 39:25]
  wire [1:0] _T_90; // @[Cat.scala 29:58]
  wire  _T_91; // @[Shift.scala 12:21]
  wire  _T_92; // @[Shift.scala 12:21]
  wire  _T_93; // @[LZD.scala 49:16]
  wire  _T_94; // @[LZD.scala 49:27]
  wire  _T_95; // @[LZD.scala 49:25]
  wire  _T_96; // @[LZD.scala 49:47]
  wire  _T_97; // @[LZD.scala 49:59]
  wire  _T_98; // @[LZD.scala 49:35]
  wire [2:0] _T_100; // @[Cat.scala 29:58]
  wire [2:0] _T_101; // @[convert.scala 21:22]
  wire [2:0] _T_102; // @[convert.scala 22:36]
  wire  _T_103; // @[Shift.scala 16:24]
  wire [1:0] _T_104; // @[Shift.scala 17:37]
  wire  _T_105; // @[Shift.scala 12:21]
  wire  _T_106; // @[Shift.scala 64:52]
  wire [2:0] _T_108; // @[Cat.scala 29:58]
  wire [2:0] _T_109; // @[Shift.scala 64:27]
  wire  _T_110; // @[Shift.scala 66:70]
  wire [1:0] _T_112; // @[Shift.scala 64:52]
  wire [2:0] _T_113; // @[Cat.scala 29:58]
  wire [2:0] _T_114; // @[Shift.scala 64:27]
  wire [2:0] _T_115; // @[Shift.scala 16:10]
  wire [1:0] _T_116; // @[convert.scala 23:34]
  wire  decB_fraction; // @[convert.scala 24:34]
  wire  _T_118; // @[convert.scala 25:26]
  wire [2:0] _T_120; // @[convert.scala 25:42]
  wire [1:0] _T_123; // @[convert.scala 26:67]
  wire [1:0] _T_124; // @[convert.scala 26:51]
  wire [5:0] _T_125; // @[Cat.scala 29:58]
  wire [4:0] _T_127; // @[convert.scala 29:56]
  wire  _T_128; // @[convert.scala 29:60]
  wire  _T_129; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_132; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_141; // @[Bitwise.scala 71:12]
  wire  _T_142; // @[PositDivisionSqrt.scala 80:40]
  wire [7:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_145; // @[PositDivisionSqrt.scala 82:31]
  wire [7:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_148; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_149; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_150; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_151; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_152; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_153; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_154; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_155; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_156; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_157; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [6:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_160; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_161; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_162; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_163; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_164; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_165; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_166; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_167; // @[PositDivisionSqrt.scala 117:30]
  wire [3:0] _T_169; // @[PositDivisionSqrt.scala 119:26]
  wire [3:0] _T_170; // @[PositDivisionSqrt.scala 118:20]
  wire [3:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [3:0] _T_171; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_173; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_174; // @[PositDivisionSqrt.scala 123:27]
  wire [2:0] _T_176; // @[PositDivisionSqrt.scala 123:52]
  wire [2:0] _T_177; // @[PositDivisionSqrt.scala 123:20]
  wire [3:0] _GEN_10; // @[PositDivisionSqrt.scala 122:64]
  wire [3:0] _T_178; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_180; // @[PositDivisionSqrt.scala 124:27]
  wire [3:0] _GEN_11; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _T_182; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _GEN_0; // @[PositDivisionSqrt.scala 116:29]
  wire [4:0] _T_183; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_185; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_186; // @[PositDivisionSqrt.scala 137:28]
  wire [7:0] _T_187; // @[PositDivisionSqrt.scala 146:22]
  wire [5:0] _T_188; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_189; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_190; // @[PositDivisionSqrt.scala 148:23]
  wire [7:0] _T_191; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_192; // @[PositDivisionSqrt.scala 149:23]
  wire [8:0] _T_193; // @[PositDivisionSqrt.scala 149:46]
  wire [7:0] _T_194; // @[PositDivisionSqrt.scala 149:56]
  wire [7:0] _T_195; // @[PositDivisionSqrt.scala 149:16]
  wire [7:0] _T_196; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_197; // @[PositDivisionSqrt.scala 150:17]
  wire [7:0] _T_198; // @[PositDivisionSqrt.scala 150:16]
  wire [7:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_200; // @[PositDivisionSqrt.scala 152:29]
  wire [7:0] _T_201; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_202; // @[PositDivisionSqrt.scala 153:29]
  wire [4:0] _T_203; // @[PositDivisionSqrt.scala 153:22]
  wire [7:0] _GEN_12; // @[PositDivisionSqrt.scala 152:93]
  wire [7:0] _T_204; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_206; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_207; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_208; // @[PositDivisionSqrt.scala 154:57]
  wire [7:0] _T_211; // @[Cat.scala 29:58]
  wire [7:0] _T_212; // @[PositDivisionSqrt.scala 154:22]
  wire [7:0] _T_213; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_215; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_216; // @[PositDivisionSqrt.scala 156:83]
  wire [3:0] _T_218; // @[Bitwise.scala 71:12]
  wire [6:0] bitMask; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  wire [6:0] _GEN_13; // @[PositDivisionSqrt.scala 156:53]
  wire [6:0] _T_219; // @[PositDivisionSqrt.scala 156:53]
  wire [7:0] _GEN_14; // @[PositDivisionSqrt.scala 155:51]
  wire [7:0] _T_220; // @[PositDivisionSqrt.scala 155:51]
  wire [5:0] _T_221; // @[PositDivisionSqrt.scala 157:53]
  wire [7:0] _GEN_15; // @[PositDivisionSqrt.scala 156:89]
  wire [7:0] _T_222; // @[PositDivisionSqrt.scala 156:89]
  wire [7:0] _T_223; // @[PositDivisionSqrt.scala 155:22]
  wire [7:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_225; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_226; // @[PositDivisionSqrt.scala 162:40]
  wire [7:0] _T_229; // @[PositDivisionSqrt.scala 163:97]
  wire [7:0] _T_231; // @[PositDivisionSqrt.scala 164:97]
  wire [7:0] _T_232; // @[PositDivisionSqrt.scala 161:92]
  wire [8:0] _T_237; // @[PositDivisionSqrt.scala 168:98]
  wire [7:0] _T_238; // @[PositDivisionSqrt.scala 168:108]
  wire [7:0] _T_240; // @[PositDivisionSqrt.scala 168:112]
  wire [7:0] _T_244; // @[PositDivisionSqrt.scala 169:112]
  wire [7:0] _T_245; // @[PositDivisionSqrt.scala 166:26]
  wire [7:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_246; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_247; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_249; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_250; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_251; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_252; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_253; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_255; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_256; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_257; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_258; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_259; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_262; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_263; // @[PositDivisionSqrt.scala 187:28]
  wire [7:0] _T_266; // @[PositDivisionSqrt.scala 188:47]
  wire [7:0] _T_267; // @[PositDivisionSqrt.scala 188:18]
  wire [5:0] _T_269; // @[PositDivisionSqrt.scala 189:18]
  wire [7:0] _GEN_16; // @[PositDivisionSqrt.scala 188:78]
  wire [7:0] _T_270; // @[PositDivisionSqrt.scala 188:78]
  wire [7:0] _GEN_17; // @[PositDivisionSqrt.scala 190:47]
  wire [7:0] _T_272; // @[PositDivisionSqrt.scala 190:47]
  wire [7:0] _T_273; // @[PositDivisionSqrt.scala 190:18]
  wire [7:0] _T_274; // @[PositDivisionSqrt.scala 189:78]
  wire [1:0] _T_276; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [7:0] _GEN_18; // @[PositDivisionSqrt.scala 197:25]
  wire [7:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire  _T_279; // @[PositDivisionSqrt.scala 200:97]
  wire  _T_280; // @[PositDivisionSqrt.scala 201:97]
  wire  realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_281; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_282; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_283; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_286; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_287; // @[Cat.scala 29:58]
  wire [2:0] _T_288; // @[PositDivisionSqrt.scala 209:63]
  wire [6:0] _GEN_19; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] _T_290; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [6:0] _T_292; // @[Mux.scala 87:16]
  wire [6:0] _T_293; // @[Mux.scala 87:16]
  wire [2:0] _T_294; // @[PositDivisionSqrt.scala 224:48]
  wire [2:0] _T_295; // @[PositDivisionSqrt.scala 224:64]
  wire [2:0] decQ_grs; // @[PositDivisionSqrt.scala 224:23]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [5:0] _GEN_20; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [5:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [1:0] _T_301; // @[convert.scala 46:61]
  wire [1:0] _T_302; // @[convert.scala 46:52]
  wire [1:0] _T_304; // @[convert.scala 46:42]
  wire [3:0] _T_305; // @[convert.scala 48:34]
  wire  _T_306; // @[convert.scala 49:36]
  wire [3:0] _T_308; // @[convert.scala 50:36]
  wire [3:0] _T_309; // @[convert.scala 50:36]
  wire [3:0] _T_310; // @[convert.scala 50:28]
  wire  _T_311; // @[convert.scala 51:31]
  wire  _T_312; // @[convert.scala 52:43]
  wire [7:0] _T_316; // @[Cat.scala 29:58]
  wire [3:0] _T_317; // @[Shift.scala 39:17]
  wire  _T_318; // @[Shift.scala 39:24]
  wire [2:0] _T_319; // @[Shift.scala 40:44]
  wire [3:0] _T_320; // @[Shift.scala 90:30]
  wire [3:0] _T_321; // @[Shift.scala 90:48]
  wire  _T_322; // @[Shift.scala 90:57]
  wire [3:0] _GEN_21; // @[Shift.scala 90:39]
  wire [3:0] _T_323; // @[Shift.scala 90:39]
  wire  _T_324; // @[Shift.scala 12:21]
  wire  _T_325; // @[Shift.scala 12:21]
  wire [3:0] _T_327; // @[Bitwise.scala 71:12]
  wire [7:0] _T_328; // @[Cat.scala 29:58]
  wire [7:0] _T_329; // @[Shift.scala 91:22]
  wire [1:0] _T_330; // @[Shift.scala 92:77]
  wire [5:0] _T_331; // @[Shift.scala 90:30]
  wire [1:0] _T_332; // @[Shift.scala 90:48]
  wire  _T_333; // @[Shift.scala 90:57]
  wire [5:0] _GEN_22; // @[Shift.scala 90:39]
  wire [5:0] _T_334; // @[Shift.scala 90:39]
  wire  _T_335; // @[Shift.scala 12:21]
  wire  _T_336; // @[Shift.scala 12:21]
  wire [1:0] _T_338; // @[Bitwise.scala 71:12]
  wire [7:0] _T_339; // @[Cat.scala 29:58]
  wire [7:0] _T_340; // @[Shift.scala 91:22]
  wire  _T_341; // @[Shift.scala 92:77]
  wire [6:0] _T_342; // @[Shift.scala 90:30]
  wire  _T_343; // @[Shift.scala 90:48]
  wire [6:0] _GEN_23; // @[Shift.scala 90:39]
  wire [6:0] _T_345; // @[Shift.scala 90:39]
  wire  _T_347; // @[Shift.scala 12:21]
  wire [7:0] _T_348; // @[Cat.scala 29:58]
  wire [7:0] _T_349; // @[Shift.scala 91:22]
  wire [7:0] _T_352; // @[Bitwise.scala 71:12]
  wire [7:0] _T_353; // @[Shift.scala 39:10]
  wire  _T_354; // @[convert.scala 55:31]
  wire  _T_355; // @[convert.scala 56:31]
  wire  _T_356; // @[convert.scala 57:31]
  wire  _T_357; // @[convert.scala 58:31]
  wire [4:0] _T_358; // @[convert.scala 59:69]
  wire  _T_359; // @[convert.scala 59:81]
  wire  _T_360; // @[convert.scala 59:50]
  wire  _T_362; // @[convert.scala 60:81]
  wire  _T_363; // @[convert.scala 61:44]
  wire  _T_364; // @[convert.scala 61:52]
  wire  _T_365; // @[convert.scala 61:36]
  wire  _T_366; // @[convert.scala 62:63]
  wire  _T_367; // @[convert.scala 62:103]
  wire  _T_368; // @[convert.scala 62:60]
  wire [4:0] _GEN_24; // @[convert.scala 63:56]
  wire [4:0] _T_371; // @[convert.scala 63:56]
  wire [5:0] _T_372; // @[Cat.scala 29:58]
  wire [5:0] _T_374; // @[Mux.scala 87:16]
  assign _T_1 = io_A[5]; // @[convert.scala 18:24]
  assign _T_2 = io_A[4]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[4:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[3:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[3:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7 != 2'h0; // @[LZD.scala 39:14]
  assign _T_9 = _T_7[1]; // @[LZD.scala 39:21]
  assign _T_10 = _T_7[0]; // @[LZD.scala 39:30]
  assign _T_11 = ~ _T_10; // @[LZD.scala 39:27]
  assign _T_12 = _T_9 | _T_11; // @[LZD.scala 39:25]
  assign _T_13 = {_T_8,_T_12}; // @[Cat.scala 29:58]
  assign _T_14 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_15 = _T_14 != 2'h0; // @[LZD.scala 39:14]
  assign _T_16 = _T_14[1]; // @[LZD.scala 39:21]
  assign _T_17 = _T_14[0]; // @[LZD.scala 39:30]
  assign _T_18 = ~ _T_17; // @[LZD.scala 39:27]
  assign _T_19 = _T_16 | _T_18; // @[LZD.scala 39:25]
  assign _T_20 = {_T_15,_T_19}; // @[Cat.scala 29:58]
  assign _T_21 = _T_13[1]; // @[Shift.scala 12:21]
  assign _T_22 = _T_20[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21 | _T_22; // @[LZD.scala 49:16]
  assign _T_24 = ~ _T_22; // @[LZD.scala 49:27]
  assign _T_25 = _T_21 | _T_24; // @[LZD.scala 49:25]
  assign _T_26 = _T_13[0:0]; // @[LZD.scala 49:47]
  assign _T_27 = _T_20[0:0]; // @[LZD.scala 49:59]
  assign _T_28 = _T_21 ? _T_26 : _T_27; // @[LZD.scala 49:35]
  assign _T_30 = {_T_23,_T_25,_T_28}; // @[Cat.scala 29:58]
  assign _T_31 = ~ _T_30; // @[convert.scala 21:22]
  assign _T_32 = io_A[2:0]; // @[convert.scala 22:36]
  assign _T_33 = _T_31 < 3'h3; // @[Shift.scala 16:24]
  assign _T_34 = _T_31[1:0]; // @[Shift.scala 17:37]
  assign _T_35 = _T_34[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_32[0:0]; // @[Shift.scala 64:52]
  assign _T_38 = {_T_36,2'h0}; // @[Cat.scala 29:58]
  assign _T_39 = _T_35 ? _T_38 : _T_32; // @[Shift.scala 64:27]
  assign _T_40 = _T_34[0:0]; // @[Shift.scala 66:70]
  assign _T_42 = _T_39[1:0]; // @[Shift.scala 64:52]
  assign _T_43 = {_T_42,1'h0}; // @[Cat.scala 29:58]
  assign _T_44 = _T_40 ? _T_43 : _T_39; // @[Shift.scala 64:27]
  assign _T_45 = _T_33 ? _T_44 : 3'h0; // @[Shift.scala 16:10]
  assign _T_46 = _T_45[2:1]; // @[convert.scala 23:34]
  assign decA_fraction = _T_45[0:0]; // @[convert.scala 24:34]
  assign _T_48 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_50 = _T_3 ? _T_31 : _T_30; // @[convert.scala 25:42]
  assign _T_53 = ~ _T_46; // @[convert.scala 26:67]
  assign _T_54 = _T_1 ? _T_53 : _T_46; // @[convert.scala 26:51]
  assign _T_55 = {_T_48,_T_50,_T_54}; // @[Cat.scala 29:58]
  assign _T_57 = io_A[4:0]; // @[convert.scala 29:56]
  assign _T_58 = _T_57 != 5'h0; // @[convert.scala 29:60]
  assign _T_59 = ~ _T_58; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_59; // @[convert.scala 29:39]
  assign _T_62 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_62 & _T_59; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_55); // @[convert.scala 32:24]
  assign _T_71 = io_B[5]; // @[convert.scala 18:24]
  assign _T_72 = io_B[4]; // @[convert.scala 18:40]
  assign _T_73 = _T_71 ^ _T_72; // @[convert.scala 18:36]
  assign _T_74 = io_B[4:1]; // @[convert.scala 19:24]
  assign _T_75 = io_B[3:0]; // @[convert.scala 19:43]
  assign _T_76 = _T_74 ^ _T_75; // @[convert.scala 19:39]
  assign _T_77 = _T_76[3:2]; // @[LZD.scala 43:32]
  assign _T_78 = _T_77 != 2'h0; // @[LZD.scala 39:14]
  assign _T_79 = _T_77[1]; // @[LZD.scala 39:21]
  assign _T_80 = _T_77[0]; // @[LZD.scala 39:30]
  assign _T_81 = ~ _T_80; // @[LZD.scala 39:27]
  assign _T_82 = _T_79 | _T_81; // @[LZD.scala 39:25]
  assign _T_83 = {_T_78,_T_82}; // @[Cat.scala 29:58]
  assign _T_84 = _T_76[1:0]; // @[LZD.scala 44:32]
  assign _T_85 = _T_84 != 2'h0; // @[LZD.scala 39:14]
  assign _T_86 = _T_84[1]; // @[LZD.scala 39:21]
  assign _T_87 = _T_84[0]; // @[LZD.scala 39:30]
  assign _T_88 = ~ _T_87; // @[LZD.scala 39:27]
  assign _T_89 = _T_86 | _T_88; // @[LZD.scala 39:25]
  assign _T_90 = {_T_85,_T_89}; // @[Cat.scala 29:58]
  assign _T_91 = _T_83[1]; // @[Shift.scala 12:21]
  assign _T_92 = _T_90[1]; // @[Shift.scala 12:21]
  assign _T_93 = _T_91 | _T_92; // @[LZD.scala 49:16]
  assign _T_94 = ~ _T_92; // @[LZD.scala 49:27]
  assign _T_95 = _T_91 | _T_94; // @[LZD.scala 49:25]
  assign _T_96 = _T_83[0:0]; // @[LZD.scala 49:47]
  assign _T_97 = _T_90[0:0]; // @[LZD.scala 49:59]
  assign _T_98 = _T_91 ? _T_96 : _T_97; // @[LZD.scala 49:35]
  assign _T_100 = {_T_93,_T_95,_T_98}; // @[Cat.scala 29:58]
  assign _T_101 = ~ _T_100; // @[convert.scala 21:22]
  assign _T_102 = io_B[2:0]; // @[convert.scala 22:36]
  assign _T_103 = _T_101 < 3'h3; // @[Shift.scala 16:24]
  assign _T_104 = _T_101[1:0]; // @[Shift.scala 17:37]
  assign _T_105 = _T_104[1]; // @[Shift.scala 12:21]
  assign _T_106 = _T_102[0:0]; // @[Shift.scala 64:52]
  assign _T_108 = {_T_106,2'h0}; // @[Cat.scala 29:58]
  assign _T_109 = _T_105 ? _T_108 : _T_102; // @[Shift.scala 64:27]
  assign _T_110 = _T_104[0:0]; // @[Shift.scala 66:70]
  assign _T_112 = _T_109[1:0]; // @[Shift.scala 64:52]
  assign _T_113 = {_T_112,1'h0}; // @[Cat.scala 29:58]
  assign _T_114 = _T_110 ? _T_113 : _T_109; // @[Shift.scala 64:27]
  assign _T_115 = _T_103 ? _T_114 : 3'h0; // @[Shift.scala 16:10]
  assign _T_116 = _T_115[2:1]; // @[convert.scala 23:34]
  assign decB_fraction = _T_115[0:0]; // @[convert.scala 24:34]
  assign _T_118 = _T_73 == 1'h0; // @[convert.scala 25:26]
  assign _T_120 = _T_73 ? _T_101 : _T_100; // @[convert.scala 25:42]
  assign _T_123 = ~ _T_116; // @[convert.scala 26:67]
  assign _T_124 = _T_71 ? _T_123 : _T_116; // @[convert.scala 26:51]
  assign _T_125 = {_T_118,_T_120,_T_124}; // @[Cat.scala 29:58]
  assign _T_127 = io_B[4:0]; // @[convert.scala 29:56]
  assign _T_128 = _T_127 != 5'h0; // @[convert.scala 29:60]
  assign _T_129 = ~ _T_128; // @[convert.scala 29:41]
  assign decB_isNaR = _T_71 & _T_129; // @[convert.scala 29:39]
  assign _T_132 = _T_71 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_132 & _T_129; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_125); // @[convert.scala 32:24]
  assign _T_141 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_142 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_141,_T_142,decA_fraction,3'h0}; // @[Cat.scala 29:58]
  assign _T_145 = ~ _T_71; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_71,_T_145,decB_fraction,5'h0}; // @[Cat.scala 29:58]
  assign _T_148 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_148 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_149 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_150 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_151 = _T_150 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_152 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_153 = decA_isZero & _T_152; // @[PositDivisionSqrt.scala 94:43]
  assign _T_154 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_155 = _T_153 & _T_154; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_156 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_157 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_156 & _T_157; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_156 & _T_62; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_160 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_160; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 3'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 3'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_161 = sigX_Z[7]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_162 = sigX_Z[5]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_161 ^ _T_162; // @[PositDivisionSqrt.scala 113:50]
  assign _T_163 = cycleNum == 3'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_163 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_164 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_165 = _T_164 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_166 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_167 = entering & _T_166; // @[PositDivisionSqrt.scala 117:30]
  assign _T_169 = io_sqrtOp ? 4'h6 : 4'h8; // @[PositDivisionSqrt.scala 119:26]
  assign _T_170 = entering_normalCase ? _T_169 : 4'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{3'd0}, _T_167}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_171 = _GEN_9 | _T_170; // @[PositDivisionSqrt.scala 117:64]
  assign _T_173 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_174 = _T_164 & _T_173; // @[PositDivisionSqrt.scala 123:27]
  assign _T_176 = cycleNum - 3'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_177 = _T_174 ? _T_176 : 3'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _GEN_10 = {{1'd0}, _T_177}; // @[PositDivisionSqrt.scala 122:64]
  assign _T_178 = _T_171 | _GEN_10; // @[PositDivisionSqrt.scala 122:64]
  assign _T_180 = _T_164 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_11 = {{3'd0}, _T_180}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_182 = _T_178 | _GEN_11; // @[PositDivisionSqrt.scala 123:64]
  assign _GEN_0 = _T_165 ? _T_182 : {{1'd0}, cycleNum}; // @[PositDivisionSqrt.scala 116:29]
  assign _T_183 = decA_scale[5:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_185 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_186 = entering_normalCase & _T_185; // @[PositDivisionSqrt.scala 137:28]
  assign _T_187 = 8'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign _T_188 = _T_187[7:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_189 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_190 = ready & _T_189; // @[PositDivisionSqrt.scala 148:23]
  assign _T_191 = _T_190 ? sigA_S : 8'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_192 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_193 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_194 = _T_193[7:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_195 = _T_192 ? _T_194 : 8'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_196 = _T_191 | _T_195; // @[PositDivisionSqrt.scala 148:66]
  assign _T_197 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_198 = _T_197 ? rem_Z : 8'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_196 | _T_198; // @[PositDivisionSqrt.scala 149:66]
  assign _T_200 = ready & _T_185; // @[PositDivisionSqrt.scala 152:29]
  assign _T_201 = _T_200 ? sigB_S : 8'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_202 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_203 = _T_202 ? 5'h10 : 5'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_12 = {{3'd0}, _T_203}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_204 = _T_201 | _GEN_12; // @[PositDivisionSqrt.scala 152:93]
  assign _T_206 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_207 = _T_197 & _T_206; // @[PositDivisionSqrt.scala 154:30]
  assign _T_208 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_211 = {signB_Z,_T_208,fractB_Z,5'h0}; // @[Cat.scala 29:58]
  assign _T_212 = _T_207 ? _T_211 : 8'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_213 = _T_204 | _T_212; // @[PositDivisionSqrt.scala 153:93]
  assign _T_215 = _T_197 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_216 = rem[7:7]; // @[PositDivisionSqrt.scala 156:83]
  assign _T_218 = _T_216 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign bitMask = {{1'd0}, _T_188}; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  assign _GEN_13 = {{3'd0}, _T_218}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_219 = bitMask & _GEN_13; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_14 = {{1'd0}, _T_219}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_220 = sigX_Z | _GEN_14; // @[PositDivisionSqrt.scala 155:51]
  assign _T_221 = bitMask[6:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_15 = {{2'd0}, _T_221}; // @[PositDivisionSqrt.scala 156:89]
  assign _T_222 = _T_220 | _GEN_15; // @[PositDivisionSqrt.scala 156:89]
  assign _T_223 = _T_215 ? _T_222 : 8'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_213 | _T_223; // @[PositDivisionSqrt.scala 154:93]
  assign _T_225 = trialTerm[7:7]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_226 = _T_216 ^ _T_225; // @[PositDivisionSqrt.scala 162:40]
  assign _T_229 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_231 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_232 = _T_226 ? _T_229 : _T_231; // @[PositDivisionSqrt.scala 161:92]
  assign _T_237 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_238 = _T_237[7:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_240 = _T_238 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_244 = _T_238 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_245 = _T_226 ? _T_240 : _T_244; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_232 : _T_245; // @[PositDivisionSqrt.scala 159:27]
  assign _T_246 = trialRem != 8'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_246 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_247 = rem != 8'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_247 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_249 = trialRem[7:7]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_250 = _T_225 ^ _T_249; // @[PositDivisionSqrt.scala 176:49]
  assign _T_251 = ~ _T_250; // @[PositDivisionSqrt.scala 176:29]
  assign _T_252 = sigX_Z[7:7]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_253 = ~ _T_252; // @[PositDivisionSqrt.scala 178:49]
  assign _T_255 = remIsZero ? _T_252 : _T_251; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_253 : _T_255; // @[Mux.scala 87:16]
  assign _T_256 = cycleNum > 3'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_257 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_258 = _T_256 & _T_257; // @[PositDivisionSqrt.scala 183:48]
  assign _T_259 = entering_normalCase | _T_258; // @[PositDivisionSqrt.scala 183:28]
  assign _T_262 = _T_197 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_263 = entering_normalCase | _T_262; // @[PositDivisionSqrt.scala 187:28]
  assign _T_266 = {newBit, 7'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_267 = _T_200 ? _T_266 : 8'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_269 = _T_202 ? 6'h20 : 6'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_16 = {{2'd0}, _T_269}; // @[PositDivisionSqrt.scala 188:78]
  assign _T_270 = _T_267 | _GEN_16; // @[PositDivisionSqrt.scala 188:78]
  assign _GEN_17 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_272 = sigX_Z | _GEN_17; // @[PositDivisionSqrt.scala 190:47]
  assign _T_273 = _T_197 ? _T_272 : 8'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_274 = _T_270 | _T_273; // @[PositDivisionSqrt.scala 189:78]
  assign _T_276 = {_T_252, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_276 : {{1'd0}, _T_252}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_18 = {{6'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_18; // @[PositDivisionSqrt.scala 197:25]
  assign _T_279 = realSigX[4]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_280 = realSigX[3]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_279 : _T_280; // @[PositDivisionSqrt.scala 198:21]
  assign _T_281 = realSigX[7]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_282 = realSigX[5]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_283 = _T_281 ^ _T_282; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_283; // @[PositDivisionSqrt.scala 205:23]
  assign notNeedSubTwo = _T_281 ^ _T_279; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_286 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_286; // @[PositDivisionSqrt.scala 208:36]
  assign _T_287 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_288 = {1'b0,$signed(_T_287)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_19 = {{4{_T_288[2]}},_T_288}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_290 = $signed(scale_Z) - $signed(_GEN_19); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_290); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-7'sh11); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(7'sh10); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[7:7]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_292 = underflow ? $signed(-7'sh11) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_293 = overflow ? $signed(7'sh10) : $signed(_T_292); // @[Mux.scala 87:16]
  assign _T_294 = realSigX[3:1]; // @[PositDivisionSqrt.scala 224:48]
  assign _T_295 = realSigX[2:0]; // @[PositDivisionSqrt.scala 224:64]
  assign decQ_grs = scaleNotChange ? _T_294 : _T_295; // @[PositDivisionSqrt.scala 224:23]
  assign outValid = cycleNum == 3'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_20 = _T_293[5:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_20); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_301 = decQ_scale[1:0]; // @[convert.scala 46:61]
  assign _T_302 = ~ _T_301; // @[convert.scala 46:52]
  assign _T_304 = decQ_sign ? _T_302 : _T_301; // @[convert.scala 46:42]
  assign _T_305 = decQ_scale[5:2]; // @[convert.scala 48:34]
  assign _T_306 = _T_305[3:3]; // @[convert.scala 49:36]
  assign _T_308 = ~ _T_305; // @[convert.scala 50:36]
  assign _T_309 = $signed(_T_308); // @[convert.scala 50:36]
  assign _T_310 = _T_306 ? $signed(_T_309) : $signed(_T_305); // @[convert.scala 50:28]
  assign _T_311 = _T_306 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_312 = ~ _T_311; // @[convert.scala 52:43]
  assign _T_316 = {_T_312,_T_311,_T_304,realFrac,decQ_grs}; // @[Cat.scala 29:58]
  assign _T_317 = $unsigned(_T_310); // @[Shift.scala 39:17]
  assign _T_318 = _T_317 < 4'h8; // @[Shift.scala 39:24]
  assign _T_319 = _T_310[2:0]; // @[Shift.scala 40:44]
  assign _T_320 = _T_316[7:4]; // @[Shift.scala 90:30]
  assign _T_321 = _T_316[3:0]; // @[Shift.scala 90:48]
  assign _T_322 = _T_321 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{3'd0}, _T_322}; // @[Shift.scala 90:39]
  assign _T_323 = _T_320 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_324 = _T_319[2]; // @[Shift.scala 12:21]
  assign _T_325 = _T_316[7]; // @[Shift.scala 12:21]
  assign _T_327 = _T_325 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_328 = {_T_327,_T_323}; // @[Cat.scala 29:58]
  assign _T_329 = _T_324 ? _T_328 : _T_316; // @[Shift.scala 91:22]
  assign _T_330 = _T_319[1:0]; // @[Shift.scala 92:77]
  assign _T_331 = _T_329[7:2]; // @[Shift.scala 90:30]
  assign _T_332 = _T_329[1:0]; // @[Shift.scala 90:48]
  assign _T_333 = _T_332 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{5'd0}, _T_333}; // @[Shift.scala 90:39]
  assign _T_334 = _T_331 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_335 = _T_330[1]; // @[Shift.scala 12:21]
  assign _T_336 = _T_329[7]; // @[Shift.scala 12:21]
  assign _T_338 = _T_336 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_339 = {_T_338,_T_334}; // @[Cat.scala 29:58]
  assign _T_340 = _T_335 ? _T_339 : _T_329; // @[Shift.scala 91:22]
  assign _T_341 = _T_330[0:0]; // @[Shift.scala 92:77]
  assign _T_342 = _T_340[7:1]; // @[Shift.scala 90:30]
  assign _T_343 = _T_340[0:0]; // @[Shift.scala 90:48]
  assign _GEN_23 = {{6'd0}, _T_343}; // @[Shift.scala 90:39]
  assign _T_345 = _T_342 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_347 = _T_340[7]; // @[Shift.scala 12:21]
  assign _T_348 = {_T_347,_T_345}; // @[Cat.scala 29:58]
  assign _T_349 = _T_341 ? _T_348 : _T_340; // @[Shift.scala 91:22]
  assign _T_352 = _T_325 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_353 = _T_318 ? _T_349 : _T_352; // @[Shift.scala 39:10]
  assign _T_354 = _T_353[3]; // @[convert.scala 55:31]
  assign _T_355 = _T_353[2]; // @[convert.scala 56:31]
  assign _T_356 = _T_353[1]; // @[convert.scala 57:31]
  assign _T_357 = _T_353[0]; // @[convert.scala 58:31]
  assign _T_358 = _T_353[7:3]; // @[convert.scala 59:69]
  assign _T_359 = _T_358 != 5'h0; // @[convert.scala 59:81]
  assign _T_360 = ~ _T_359; // @[convert.scala 59:50]
  assign _T_362 = _T_358 == 5'h1f; // @[convert.scala 60:81]
  assign _T_363 = _T_354 | _T_356; // @[convert.scala 61:44]
  assign _T_364 = _T_363 | _T_357; // @[convert.scala 61:52]
  assign _T_365 = _T_355 & _T_364; // @[convert.scala 61:36]
  assign _T_366 = ~ _T_362; // @[convert.scala 62:63]
  assign _T_367 = _T_366 & _T_365; // @[convert.scala 62:103]
  assign _T_368 = _T_360 | _T_367; // @[convert.scala 62:60]
  assign _GEN_24 = {{4'd0}, _T_368}; // @[convert.scala 63:56]
  assign _T_371 = _T_358 + _GEN_24; // @[convert.scala 63:56]
  assign _T_372 = {decQ_sign,_T_371}; // @[Cat.scala 29:58]
  assign _T_374 = isZero_Z ? 6'h0 : _T_372; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 3'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_206; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 6'h20 : _T_374; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 3'h0;
    end else begin
      cycleNum <= _GEN_0[2:0];
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_149;
      end else begin
        isNaR_Z <= _T_151;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_155;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_183[4]}},_T_183};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_186) begin
      signB_Z <= _T_71;
    end
    if (_T_186) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_259) begin
      if (ready) begin
        if (_T_226) begin
          rem_Z <= _T_229;
        end else begin
          rem_Z <= _T_231;
        end
      end else begin
        if (_T_226) begin
          rem_Z <= _T_240;
        end else begin
          rem_Z <= _T_244;
        end
      end
    end
    if (_T_263) begin
      sigX_Z <= _T_274;
    end
  end
endmodule
