module Shifter7_7(
  input        clock,
  input        reset,
  input  [6:0] io_in,
  input  [6:0] io_shiftamt,
  output [6:0] io_shiftout
);
  wire  _T; // @[Shift.scala 39:24]
  wire [2:0] _T_1; // @[Shift.scala 40:44]
  wire [2:0] _T_2; // @[Shift.scala 90:30]
  wire [3:0] _T_3; // @[Shift.scala 90:48]
  wire  _T_4; // @[Shift.scala 90:57]
  wire [2:0] _GEN_0; // @[Shift.scala 90:39]
  wire [2:0] _T_5; // @[Shift.scala 90:39]
  wire  _T_6; // @[Shift.scala 12:21]
  wire  _T_7; // @[Shift.scala 12:21]
  wire [3:0] _T_9; // @[Bitwise.scala 71:12]
  wire [6:0] _T_10; // @[Cat.scala 29:58]
  wire [6:0] _T_11; // @[Shift.scala 91:22]
  wire [1:0] _T_12; // @[Shift.scala 92:77]
  wire [4:0] _T_13; // @[Shift.scala 90:30]
  wire [1:0] _T_14; // @[Shift.scala 90:48]
  wire  _T_15; // @[Shift.scala 90:57]
  wire [4:0] _GEN_1; // @[Shift.scala 90:39]
  wire [4:0] _T_16; // @[Shift.scala 90:39]
  wire  _T_17; // @[Shift.scala 12:21]
  wire  _T_18; // @[Shift.scala 12:21]
  wire [1:0] _T_20; // @[Bitwise.scala 71:12]
  wire [6:0] _T_21; // @[Cat.scala 29:58]
  wire [6:0] _T_22; // @[Shift.scala 91:22]
  wire  _T_23; // @[Shift.scala 92:77]
  wire [5:0] _T_24; // @[Shift.scala 90:30]
  wire  _T_25; // @[Shift.scala 90:48]
  wire [5:0] _GEN_2; // @[Shift.scala 90:39]
  wire [5:0] _T_27; // @[Shift.scala 90:39]
  wire  _T_29; // @[Shift.scala 12:21]
  wire [6:0] _T_30; // @[Cat.scala 29:58]
  wire [6:0] _T_31; // @[Shift.scala 91:22]
  wire [6:0] _T_34; // @[Bitwise.scala 71:12]
  assign _T = io_shiftamt < 7'h7; // @[Shift.scala 39:24]
  assign _T_1 = io_shiftamt[2:0]; // @[Shift.scala 40:44]
  assign _T_2 = io_in[6:4]; // @[Shift.scala 90:30]
  assign _T_3 = io_in[3:0]; // @[Shift.scala 90:48]
  assign _T_4 = _T_3 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{2'd0}, _T_4}; // @[Shift.scala 90:39]
  assign _T_5 = _T_2 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_6 = _T_1[2]; // @[Shift.scala 12:21]
  assign _T_7 = io_in[6]; // @[Shift.scala 12:21]
  assign _T_9 = _T_7 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_10 = {_T_9,_T_5}; // @[Cat.scala 29:58]
  assign _T_11 = _T_6 ? _T_10 : io_in; // @[Shift.scala 91:22]
  assign _T_12 = _T_1[1:0]; // @[Shift.scala 92:77]
  assign _T_13 = _T_11[6:2]; // @[Shift.scala 90:30]
  assign _T_14 = _T_11[1:0]; // @[Shift.scala 90:48]
  assign _T_15 = _T_14 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{4'd0}, _T_15}; // @[Shift.scala 90:39]
  assign _T_16 = _T_13 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_17 = _T_12[1]; // @[Shift.scala 12:21]
  assign _T_18 = _T_11[6]; // @[Shift.scala 12:21]
  assign _T_20 = _T_18 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_21 = {_T_20,_T_16}; // @[Cat.scala 29:58]
  assign _T_22 = _T_17 ? _T_21 : _T_11; // @[Shift.scala 91:22]
  assign _T_23 = _T_12[0:0]; // @[Shift.scala 92:77]
  assign _T_24 = _T_22[6:1]; // @[Shift.scala 90:30]
  assign _T_25 = _T_22[0:0]; // @[Shift.scala 90:48]
  assign _GEN_2 = {{5'd0}, _T_25}; // @[Shift.scala 90:39]
  assign _T_27 = _T_24 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_29 = _T_22[6]; // @[Shift.scala 12:21]
  assign _T_30 = {_T_29,_T_27}; // @[Cat.scala 29:58]
  assign _T_31 = _T_23 ? _T_30 : _T_22; // @[Shift.scala 91:22]
  assign _T_34 = _T_7 ? 7'h7f : 7'h0; // @[Bitwise.scala 71:12]
  assign io_shiftout = _T ? _T_31 : _T_34; // @[Shif.scala 16:15]
endmodule
