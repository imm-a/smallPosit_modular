module Sig_op8_0(
  input        clock,
  input        reset,
  input  [7:0] io_A,
  input  [7:0] io_B,
  output       io_greaterSign,
  output       io_smallerSign,
  output [3:0] io_greaterExp,
  output [6:0] io_greaterSig,
  output [9:0] io_smallerSig,
  output       io_AisNar,
  output       io_BisNar,
  output       io_AisZero,
  output       io_BisZero
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [5:0] _T_4; // @[convert.scala 19:24]
  wire [5:0] _T_5; // @[convert.scala 19:43]
  wire [5:0] _T_6; // @[convert.scala 19:39]
  wire [3:0] _T_7; // @[LZD.scala 43:32]
  wire [1:0] _T_8; // @[LZD.scala 43:32]
  wire  _T_9; // @[LZD.scala 39:14]
  wire  _T_10; // @[LZD.scala 39:21]
  wire  _T_11; // @[LZD.scala 39:30]
  wire  _T_12; // @[LZD.scala 39:27]
  wire  _T_13; // @[LZD.scala 39:25]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [1:0] _T_15; // @[LZD.scala 44:32]
  wire  _T_16; // @[LZD.scala 39:14]
  wire  _T_17; // @[LZD.scala 39:21]
  wire  _T_18; // @[LZD.scala 39:30]
  wire  _T_19; // @[LZD.scala 39:27]
  wire  _T_20; // @[LZD.scala 39:25]
  wire [1:0] _T_21; // @[Cat.scala 29:58]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[LZD.scala 49:16]
  wire  _T_25; // @[LZD.scala 49:27]
  wire  _T_26; // @[LZD.scala 49:25]
  wire  _T_27; // @[LZD.scala 49:47]
  wire  _T_28; // @[LZD.scala 49:59]
  wire  _T_29; // @[LZD.scala 49:35]
  wire [2:0] _T_31; // @[Cat.scala 29:58]
  wire [1:0] _T_32; // @[LZD.scala 44:32]
  wire  _T_33; // @[LZD.scala 39:14]
  wire  _T_34; // @[LZD.scala 39:21]
  wire  _T_35; // @[LZD.scala 39:30]
  wire  _T_36; // @[LZD.scala 39:27]
  wire  _T_37; // @[LZD.scala 39:25]
  wire [1:0] _T_38; // @[Cat.scala 29:58]
  wire  _T_39; // @[Shift.scala 12:21]
  wire [1:0] _T_41; // @[LZD.scala 55:32]
  wire [1:0] _T_42; // @[LZD.scala 55:20]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire [2:0] _T_44; // @[convert.scala 21:22]
  wire [4:0] _T_45; // @[convert.scala 22:36]
  wire  _T_46; // @[Shift.scala 16:24]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 64:52]
  wire [4:0] _T_51; // @[Cat.scala 29:58]
  wire [4:0] _T_52; // @[Shift.scala 64:27]
  wire [1:0] _T_53; // @[Shift.scala 66:70]
  wire  _T_54; // @[Shift.scala 12:21]
  wire [2:0] _T_55; // @[Shift.scala 64:52]
  wire [4:0] _T_57; // @[Cat.scala 29:58]
  wire [4:0] _T_58; // @[Shift.scala 64:27]
  wire  _T_59; // @[Shift.scala 66:70]
  wire [3:0] _T_61; // @[Shift.scala 64:52]
  wire [4:0] _T_62; // @[Cat.scala 29:58]
  wire [4:0] _T_63; // @[Shift.scala 64:27]
  wire [4:0] decA_fraction; // @[Shift.scala 16:10]
  wire  _T_67; // @[convert.scala 25:26]
  wire [2:0] _T_69; // @[convert.scala 25:42]
  wire [3:0] _T_70; // @[Cat.scala 29:58]
  wire [6:0] _T_72; // @[convert.scala 29:56]
  wire  _T_73; // @[convert.scala 29:60]
  wire  _T_74; // @[convert.scala 29:41]
  wire  _T_77; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [3:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_86; // @[convert.scala 18:24]
  wire  _T_87; // @[convert.scala 18:40]
  wire  _T_88; // @[convert.scala 18:36]
  wire [5:0] _T_89; // @[convert.scala 19:24]
  wire [5:0] _T_90; // @[convert.scala 19:43]
  wire [5:0] _T_91; // @[convert.scala 19:39]
  wire [3:0] _T_92; // @[LZD.scala 43:32]
  wire [1:0] _T_93; // @[LZD.scala 43:32]
  wire  _T_94; // @[LZD.scala 39:14]
  wire  _T_95; // @[LZD.scala 39:21]
  wire  _T_96; // @[LZD.scala 39:30]
  wire  _T_97; // @[LZD.scala 39:27]
  wire  _T_98; // @[LZD.scala 39:25]
  wire [1:0] _T_99; // @[Cat.scala 29:58]
  wire [1:0] _T_100; // @[LZD.scala 44:32]
  wire  _T_101; // @[LZD.scala 39:14]
  wire  _T_102; // @[LZD.scala 39:21]
  wire  _T_103; // @[LZD.scala 39:30]
  wire  _T_104; // @[LZD.scala 39:27]
  wire  _T_105; // @[LZD.scala 39:25]
  wire [1:0] _T_106; // @[Cat.scala 29:58]
  wire  _T_107; // @[Shift.scala 12:21]
  wire  _T_108; // @[Shift.scala 12:21]
  wire  _T_109; // @[LZD.scala 49:16]
  wire  _T_110; // @[LZD.scala 49:27]
  wire  _T_111; // @[LZD.scala 49:25]
  wire  _T_112; // @[LZD.scala 49:47]
  wire  _T_113; // @[LZD.scala 49:59]
  wire  _T_114; // @[LZD.scala 49:35]
  wire [2:0] _T_116; // @[Cat.scala 29:58]
  wire [1:0] _T_117; // @[LZD.scala 44:32]
  wire  _T_118; // @[LZD.scala 39:14]
  wire  _T_119; // @[LZD.scala 39:21]
  wire  _T_120; // @[LZD.scala 39:30]
  wire  _T_121; // @[LZD.scala 39:27]
  wire  _T_122; // @[LZD.scala 39:25]
  wire [1:0] _T_123; // @[Cat.scala 29:58]
  wire  _T_124; // @[Shift.scala 12:21]
  wire [1:0] _T_126; // @[LZD.scala 55:32]
  wire [1:0] _T_127; // @[LZD.scala 55:20]
  wire [2:0] _T_128; // @[Cat.scala 29:58]
  wire [2:0] _T_129; // @[convert.scala 21:22]
  wire [4:0] _T_130; // @[convert.scala 22:36]
  wire  _T_131; // @[Shift.scala 16:24]
  wire  _T_133; // @[Shift.scala 12:21]
  wire  _T_134; // @[Shift.scala 64:52]
  wire [4:0] _T_136; // @[Cat.scala 29:58]
  wire [4:0] _T_137; // @[Shift.scala 64:27]
  wire [1:0] _T_138; // @[Shift.scala 66:70]
  wire  _T_139; // @[Shift.scala 12:21]
  wire [2:0] _T_140; // @[Shift.scala 64:52]
  wire [4:0] _T_142; // @[Cat.scala 29:58]
  wire [4:0] _T_143; // @[Shift.scala 64:27]
  wire  _T_144; // @[Shift.scala 66:70]
  wire [3:0] _T_146; // @[Shift.scala 64:52]
  wire [4:0] _T_147; // @[Cat.scala 29:58]
  wire [4:0] _T_148; // @[Shift.scala 64:27]
  wire [4:0] decB_fraction; // @[Shift.scala 16:10]
  wire  _T_152; // @[convert.scala 25:26]
  wire [2:0] _T_154; // @[convert.scala 25:42]
  wire [3:0] _T_155; // @[Cat.scala 29:58]
  wire [6:0] _T_157; // @[convert.scala 29:56]
  wire  _T_158; // @[convert.scala 29:60]
  wire  _T_159; // @[convert.scala 29:41]
  wire  _T_162; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [3:0] decB_scale; // @[convert.scala 32:24]
  wire  aGTb; // @[Sig_op.scala 38:32]
  wire [3:0] smallerExp; // @[Sig_op.scala 42:24]
  wire [4:0] greaterFrac; // @[Sig_op.scala 43:24]
  wire [4:0] smallerFrac; // @[Sig_op.scala 44:24]
  wire  smallerZero; // @[Sig_op.scala 45:24]
  wire [3:0] _T_174; // @[Sig_op.scala 46:35]
  wire [3:0] scale_diff; // @[Sig_op.scala 46:35]
  wire  _T_175; // @[Sig_op.scala 51:53]
  wire  _T_176; // @[Sig_op.scala 51:36]
  wire [9:0] _T_179; // @[Cat.scala 29:58]
  wire [3:0] _T_180; // @[Sig_op.scala 51:124]
  wire  _T_181; // @[Shift.scala 39:24]
  wire [1:0] _T_183; // @[Shift.scala 90:30]
  wire [7:0] _T_184; // @[Shift.scala 90:48]
  wire  _T_185; // @[Shift.scala 90:57]
  wire [1:0] _GEN_0; // @[Shift.scala 90:39]
  wire [1:0] _T_186; // @[Shift.scala 90:39]
  wire  _T_187; // @[Shift.scala 12:21]
  wire  _T_188; // @[Shift.scala 12:21]
  wire [7:0] _T_190; // @[Bitwise.scala 71:12]
  wire [9:0] _T_191; // @[Cat.scala 29:58]
  wire [9:0] _T_192; // @[Shift.scala 91:22]
  wire [2:0] _T_193; // @[Shift.scala 92:77]
  wire [5:0] _T_194; // @[Shift.scala 90:30]
  wire [3:0] _T_195; // @[Shift.scala 90:48]
  wire  _T_196; // @[Shift.scala 90:57]
  wire [5:0] _GEN_1; // @[Shift.scala 90:39]
  wire [5:0] _T_197; // @[Shift.scala 90:39]
  wire  _T_198; // @[Shift.scala 12:21]
  wire  _T_199; // @[Shift.scala 12:21]
  wire [3:0] _T_201; // @[Bitwise.scala 71:12]
  wire [9:0] _T_202; // @[Cat.scala 29:58]
  wire [9:0] _T_203; // @[Shift.scala 91:22]
  wire [1:0] _T_204; // @[Shift.scala 92:77]
  wire [7:0] _T_205; // @[Shift.scala 90:30]
  wire [1:0] _T_206; // @[Shift.scala 90:48]
  wire  _T_207; // @[Shift.scala 90:57]
  wire [7:0] _GEN_2; // @[Shift.scala 90:39]
  wire [7:0] _T_208; // @[Shift.scala 90:39]
  wire  _T_209; // @[Shift.scala 12:21]
  wire  _T_210; // @[Shift.scala 12:21]
  wire [1:0] _T_212; // @[Bitwise.scala 71:12]
  wire [9:0] _T_213; // @[Cat.scala 29:58]
  wire [9:0] _T_214; // @[Shift.scala 91:22]
  wire  _T_215; // @[Shift.scala 92:77]
  wire [8:0] _T_216; // @[Shift.scala 90:30]
  wire  _T_217; // @[Shift.scala 90:48]
  wire [8:0] _GEN_3; // @[Shift.scala 90:39]
  wire [8:0] _T_219; // @[Shift.scala 90:39]
  wire  _T_221; // @[Shift.scala 12:21]
  wire [9:0] _T_222; // @[Cat.scala 29:58]
  wire [9:0] _T_223; // @[Shift.scala 91:22]
  wire [9:0] _T_226; // @[Bitwise.scala 71:12]
  wire  _T_227; // @[Sig_op.scala 57:40]
  wire [1:0] _T_228; // @[Cat.scala 29:58]
  assign _T_1 = io_A[7]; // @[convert.scala 18:24]
  assign _T_2 = io_A[6]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[6:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[5:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[5:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[3:2]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8 != 2'h0; // @[LZD.scala 39:14]
  assign _T_10 = _T_8[1]; // @[LZD.scala 39:21]
  assign _T_11 = _T_8[0]; // @[LZD.scala 39:30]
  assign _T_12 = ~ _T_11; // @[LZD.scala 39:27]
  assign _T_13 = _T_10 | _T_12; // @[LZD.scala 39:25]
  assign _T_14 = {_T_9,_T_13}; // @[Cat.scala 29:58]
  assign _T_15 = _T_7[1:0]; // @[LZD.scala 44:32]
  assign _T_16 = _T_15 != 2'h0; // @[LZD.scala 39:14]
  assign _T_17 = _T_15[1]; // @[LZD.scala 39:21]
  assign _T_18 = _T_15[0]; // @[LZD.scala 39:30]
  assign _T_19 = ~ _T_18; // @[LZD.scala 39:27]
  assign _T_20 = _T_17 | _T_19; // @[LZD.scala 39:25]
  assign _T_21 = {_T_16,_T_20}; // @[Cat.scala 29:58]
  assign _T_22 = _T_14[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22 | _T_23; // @[LZD.scala 49:16]
  assign _T_25 = ~ _T_23; // @[LZD.scala 49:27]
  assign _T_26 = _T_22 | _T_25; // @[LZD.scala 49:25]
  assign _T_27 = _T_14[0:0]; // @[LZD.scala 49:47]
  assign _T_28 = _T_21[0:0]; // @[LZD.scala 49:59]
  assign _T_29 = _T_22 ? _T_27 : _T_28; // @[LZD.scala 49:35]
  assign _T_31 = {_T_24,_T_26,_T_29}; // @[Cat.scala 29:58]
  assign _T_32 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_33 = _T_32 != 2'h0; // @[LZD.scala 39:14]
  assign _T_34 = _T_32[1]; // @[LZD.scala 39:21]
  assign _T_35 = _T_32[0]; // @[LZD.scala 39:30]
  assign _T_36 = ~ _T_35; // @[LZD.scala 39:27]
  assign _T_37 = _T_34 | _T_36; // @[LZD.scala 39:25]
  assign _T_38 = {_T_33,_T_37}; // @[Cat.scala 29:58]
  assign _T_39 = _T_31[2]; // @[Shift.scala 12:21]
  assign _T_41 = _T_31[1:0]; // @[LZD.scala 55:32]
  assign _T_42 = _T_39 ? _T_41 : _T_38; // @[LZD.scala 55:20]
  assign _T_43 = {_T_39,_T_42}; // @[Cat.scala 29:58]
  assign _T_44 = ~ _T_43; // @[convert.scala 21:22]
  assign _T_45 = io_A[4:0]; // @[convert.scala 22:36]
  assign _T_46 = _T_44 < 3'h5; // @[Shift.scala 16:24]
  assign _T_48 = _T_44[2]; // @[Shift.scala 12:21]
  assign _T_49 = _T_45[0:0]; // @[Shift.scala 64:52]
  assign _T_51 = {_T_49,4'h0}; // @[Cat.scala 29:58]
  assign _T_52 = _T_48 ? _T_51 : _T_45; // @[Shift.scala 64:27]
  assign _T_53 = _T_44[1:0]; // @[Shift.scala 66:70]
  assign _T_54 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_55 = _T_52[2:0]; // @[Shift.scala 64:52]
  assign _T_57 = {_T_55,2'h0}; // @[Cat.scala 29:58]
  assign _T_58 = _T_54 ? _T_57 : _T_52; // @[Shift.scala 64:27]
  assign _T_59 = _T_53[0:0]; // @[Shift.scala 66:70]
  assign _T_61 = _T_58[3:0]; // @[Shift.scala 64:52]
  assign _T_62 = {_T_61,1'h0}; // @[Cat.scala 29:58]
  assign _T_63 = _T_59 ? _T_62 : _T_58; // @[Shift.scala 64:27]
  assign decA_fraction = _T_46 ? _T_63 : 5'h0; // @[Shift.scala 16:10]
  assign _T_67 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_69 = _T_3 ? _T_44 : _T_43; // @[convert.scala 25:42]
  assign _T_70 = {_T_67,_T_69}; // @[Cat.scala 29:58]
  assign _T_72 = io_A[6:0]; // @[convert.scala 29:56]
  assign _T_73 = _T_72 != 7'h0; // @[convert.scala 29:60]
  assign _T_74 = ~ _T_73; // @[convert.scala 29:41]
  assign _T_77 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_77 & _T_74; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_70); // @[convert.scala 32:24]
  assign _T_86 = io_B[7]; // @[convert.scala 18:24]
  assign _T_87 = io_B[6]; // @[convert.scala 18:40]
  assign _T_88 = _T_86 ^ _T_87; // @[convert.scala 18:36]
  assign _T_89 = io_B[6:1]; // @[convert.scala 19:24]
  assign _T_90 = io_B[5:0]; // @[convert.scala 19:43]
  assign _T_91 = _T_89 ^ _T_90; // @[convert.scala 19:39]
  assign _T_92 = _T_91[5:2]; // @[LZD.scala 43:32]
  assign _T_93 = _T_92[3:2]; // @[LZD.scala 43:32]
  assign _T_94 = _T_93 != 2'h0; // @[LZD.scala 39:14]
  assign _T_95 = _T_93[1]; // @[LZD.scala 39:21]
  assign _T_96 = _T_93[0]; // @[LZD.scala 39:30]
  assign _T_97 = ~ _T_96; // @[LZD.scala 39:27]
  assign _T_98 = _T_95 | _T_97; // @[LZD.scala 39:25]
  assign _T_99 = {_T_94,_T_98}; // @[Cat.scala 29:58]
  assign _T_100 = _T_92[1:0]; // @[LZD.scala 44:32]
  assign _T_101 = _T_100 != 2'h0; // @[LZD.scala 39:14]
  assign _T_102 = _T_100[1]; // @[LZD.scala 39:21]
  assign _T_103 = _T_100[0]; // @[LZD.scala 39:30]
  assign _T_104 = ~ _T_103; // @[LZD.scala 39:27]
  assign _T_105 = _T_102 | _T_104; // @[LZD.scala 39:25]
  assign _T_106 = {_T_101,_T_105}; // @[Cat.scala 29:58]
  assign _T_107 = _T_99[1]; // @[Shift.scala 12:21]
  assign _T_108 = _T_106[1]; // @[Shift.scala 12:21]
  assign _T_109 = _T_107 | _T_108; // @[LZD.scala 49:16]
  assign _T_110 = ~ _T_108; // @[LZD.scala 49:27]
  assign _T_111 = _T_107 | _T_110; // @[LZD.scala 49:25]
  assign _T_112 = _T_99[0:0]; // @[LZD.scala 49:47]
  assign _T_113 = _T_106[0:0]; // @[LZD.scala 49:59]
  assign _T_114 = _T_107 ? _T_112 : _T_113; // @[LZD.scala 49:35]
  assign _T_116 = {_T_109,_T_111,_T_114}; // @[Cat.scala 29:58]
  assign _T_117 = _T_91[1:0]; // @[LZD.scala 44:32]
  assign _T_118 = _T_117 != 2'h0; // @[LZD.scala 39:14]
  assign _T_119 = _T_117[1]; // @[LZD.scala 39:21]
  assign _T_120 = _T_117[0]; // @[LZD.scala 39:30]
  assign _T_121 = ~ _T_120; // @[LZD.scala 39:27]
  assign _T_122 = _T_119 | _T_121; // @[LZD.scala 39:25]
  assign _T_123 = {_T_118,_T_122}; // @[Cat.scala 29:58]
  assign _T_124 = _T_116[2]; // @[Shift.scala 12:21]
  assign _T_126 = _T_116[1:0]; // @[LZD.scala 55:32]
  assign _T_127 = _T_124 ? _T_126 : _T_123; // @[LZD.scala 55:20]
  assign _T_128 = {_T_124,_T_127}; // @[Cat.scala 29:58]
  assign _T_129 = ~ _T_128; // @[convert.scala 21:22]
  assign _T_130 = io_B[4:0]; // @[convert.scala 22:36]
  assign _T_131 = _T_129 < 3'h5; // @[Shift.scala 16:24]
  assign _T_133 = _T_129[2]; // @[Shift.scala 12:21]
  assign _T_134 = _T_130[0:0]; // @[Shift.scala 64:52]
  assign _T_136 = {_T_134,4'h0}; // @[Cat.scala 29:58]
  assign _T_137 = _T_133 ? _T_136 : _T_130; // @[Shift.scala 64:27]
  assign _T_138 = _T_129[1:0]; // @[Shift.scala 66:70]
  assign _T_139 = _T_138[1]; // @[Shift.scala 12:21]
  assign _T_140 = _T_137[2:0]; // @[Shift.scala 64:52]
  assign _T_142 = {_T_140,2'h0}; // @[Cat.scala 29:58]
  assign _T_143 = _T_139 ? _T_142 : _T_137; // @[Shift.scala 64:27]
  assign _T_144 = _T_138[0:0]; // @[Shift.scala 66:70]
  assign _T_146 = _T_143[3:0]; // @[Shift.scala 64:52]
  assign _T_147 = {_T_146,1'h0}; // @[Cat.scala 29:58]
  assign _T_148 = _T_144 ? _T_147 : _T_143; // @[Shift.scala 64:27]
  assign decB_fraction = _T_131 ? _T_148 : 5'h0; // @[Shift.scala 16:10]
  assign _T_152 = _T_88 == 1'h0; // @[convert.scala 25:26]
  assign _T_154 = _T_88 ? _T_129 : _T_128; // @[convert.scala 25:42]
  assign _T_155 = {_T_152,_T_154}; // @[Cat.scala 29:58]
  assign _T_157 = io_B[6:0]; // @[convert.scala 29:56]
  assign _T_158 = _T_157 != 7'h0; // @[convert.scala 29:60]
  assign _T_159 = ~ _T_158; // @[convert.scala 29:41]
  assign _T_162 = _T_86 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_162 & _T_159; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_155); // @[convert.scala 32:24]
  assign aGTb = $signed(decA_scale) > $signed(decB_scale); // @[Sig_op.scala 38:32]
  assign smallerExp = aGTb ? $signed(decB_scale) : $signed(decA_scale); // @[Sig_op.scala 42:24]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[Sig_op.scala 43:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[Sig_op.scala 44:24]
  assign smallerZero = aGTb ? decB_isZero : decA_isZero; // @[Sig_op.scala 45:24]
  assign _T_174 = $signed(io_greaterExp) - $signed(smallerExp); // @[Sig_op.scala 46:35]
  assign scale_diff = $signed(_T_174); // @[Sig_op.scala 46:35]
  assign _T_175 = io_smallerSign | smallerZero; // @[Sig_op.scala 51:53]
  assign _T_176 = ~ _T_175; // @[Sig_op.scala 51:36]
  assign _T_179 = {io_smallerSign,_T_176,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_180 = $unsigned(scale_diff); // @[Sig_op.scala 51:124]
  assign _T_181 = _T_180 < 4'ha; // @[Shift.scala 39:24]
  assign _T_183 = _T_179[9:8]; // @[Shift.scala 90:30]
  assign _T_184 = _T_179[7:0]; // @[Shift.scala 90:48]
  assign _T_185 = _T_184 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{1'd0}, _T_185}; // @[Shift.scala 90:39]
  assign _T_186 = _T_183 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_187 = _T_180[3]; // @[Shift.scala 12:21]
  assign _T_188 = _T_179[9]; // @[Shift.scala 12:21]
  assign _T_190 = _T_188 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_191 = {_T_190,_T_186}; // @[Cat.scala 29:58]
  assign _T_192 = _T_187 ? _T_191 : _T_179; // @[Shift.scala 91:22]
  assign _T_193 = _T_180[2:0]; // @[Shift.scala 92:77]
  assign _T_194 = _T_192[9:4]; // @[Shift.scala 90:30]
  assign _T_195 = _T_192[3:0]; // @[Shift.scala 90:48]
  assign _T_196 = _T_195 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{5'd0}, _T_196}; // @[Shift.scala 90:39]
  assign _T_197 = _T_194 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_198 = _T_193[2]; // @[Shift.scala 12:21]
  assign _T_199 = _T_192[9]; // @[Shift.scala 12:21]
  assign _T_201 = _T_199 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_202 = {_T_201,_T_197}; // @[Cat.scala 29:58]
  assign _T_203 = _T_198 ? _T_202 : _T_192; // @[Shift.scala 91:22]
  assign _T_204 = _T_193[1:0]; // @[Shift.scala 92:77]
  assign _T_205 = _T_203[9:2]; // @[Shift.scala 90:30]
  assign _T_206 = _T_203[1:0]; // @[Shift.scala 90:48]
  assign _T_207 = _T_206 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{7'd0}, _T_207}; // @[Shift.scala 90:39]
  assign _T_208 = _T_205 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_209 = _T_204[1]; // @[Shift.scala 12:21]
  assign _T_210 = _T_203[9]; // @[Shift.scala 12:21]
  assign _T_212 = _T_210 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_213 = {_T_212,_T_208}; // @[Cat.scala 29:58]
  assign _T_214 = _T_209 ? _T_213 : _T_203; // @[Shift.scala 91:22]
  assign _T_215 = _T_204[0:0]; // @[Shift.scala 92:77]
  assign _T_216 = _T_214[9:1]; // @[Shift.scala 90:30]
  assign _T_217 = _T_214[0:0]; // @[Shift.scala 90:48]
  assign _GEN_3 = {{8'd0}, _T_217}; // @[Shift.scala 90:39]
  assign _T_219 = _T_216 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_221 = _T_214[9]; // @[Shift.scala 12:21]
  assign _T_222 = {_T_221,_T_219}; // @[Cat.scala 29:58]
  assign _T_223 = _T_215 ? _T_222 : _T_214; // @[Shift.scala 91:22]
  assign _T_226 = _T_188 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_227 = ~ io_greaterSign; // @[Sig_op.scala 57:40]
  assign _T_228 = {io_greaterSign,_T_227}; // @[Cat.scala 29:58]
  assign io_greaterSign = aGTb ? _T_1 : _T_86; // @[Sig_op.scala 39:18]
  assign io_smallerSign = aGTb ? _T_86 : _T_1; // @[Sig_op.scala 40:18]
  assign io_greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[Sig_op.scala 41:18]
  assign io_greaterSig = {_T_228,greaterFrac}; // @[Sig_op.scala 57:17]
  assign io_smallerSig = _T_181 ? _T_223 : _T_226; // @[Sig_op.scala 52:17]
  assign io_AisNar = _T_1 & _T_74; // @[Sig_op.scala 47:13]
  assign io_BisNar = _T_86 & _T_159; // @[Sig_op.scala 48:13]
  assign io_AisZero = _T_77 & _T_74; // @[Sig_op.scala 49:14]
  assign io_BisZero = _T_162 & _T_159; // @[Sig_op.scala 50:14]
endmodule
