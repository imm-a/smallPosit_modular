module QuireToPosit14_8_1(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [63:0] io_quireIn,
  output [7:0]  io_positOut,
  output        io_outValid
);
  wire [62:0] _T; // @[QuireToPosit.scala 47:43]
  wire  _T_1; // @[QuireToPosit.scala 47:47]
  wire  tailIsZero; // @[QuireToPosit.scala 47:27]
  wire  _T_2; // @[QuireToPosit.scala 49:45]
  wire  outRawFloat_isNaR; // @[QuireToPosit.scala 49:49]
  wire  _T_5; // @[QuireToPosit.scala 50:31]
  wire  outRawFloat_isZero; // @[QuireToPosit.scala 50:51]
  wire [62:0] _T_8; // @[QuireToPosit.scala 58:41]
  wire [62:0] _T_9; // @[QuireToPosit.scala 58:68]
  wire [62:0] quireXOR; // @[QuireToPosit.scala 58:56]
  wire [31:0] _T_10; // @[LZD.scala 43:32]
  wire [15:0] _T_11; // @[LZD.scala 43:32]
  wire [7:0] _T_12; // @[LZD.scala 43:32]
  wire [3:0] _T_13; // @[LZD.scala 43:32]
  wire [1:0] _T_14; // @[LZD.scala 43:32]
  wire  _T_15; // @[LZD.scala 39:14]
  wire  _T_16; // @[LZD.scala 39:21]
  wire  _T_17; // @[LZD.scala 39:30]
  wire  _T_18; // @[LZD.scala 39:27]
  wire  _T_19; // @[LZD.scala 39:25]
  wire [1:0] _T_20; // @[Cat.scala 29:58]
  wire [1:0] _T_21; // @[LZD.scala 44:32]
  wire  _T_22; // @[LZD.scala 39:14]
  wire  _T_23; // @[LZD.scala 39:21]
  wire  _T_24; // @[LZD.scala 39:30]
  wire  _T_25; // @[LZD.scala 39:27]
  wire  _T_26; // @[LZD.scala 39:25]
  wire [1:0] _T_27; // @[Cat.scala 29:58]
  wire  _T_28; // @[Shift.scala 12:21]
  wire  _T_29; // @[Shift.scala 12:21]
  wire  _T_30; // @[LZD.scala 49:16]
  wire  _T_31; // @[LZD.scala 49:27]
  wire  _T_32; // @[LZD.scala 49:25]
  wire  _T_33; // @[LZD.scala 49:47]
  wire  _T_34; // @[LZD.scala 49:59]
  wire  _T_35; // @[LZD.scala 49:35]
  wire [2:0] _T_37; // @[Cat.scala 29:58]
  wire [3:0] _T_38; // @[LZD.scala 44:32]
  wire [1:0] _T_39; // @[LZD.scala 43:32]
  wire  _T_40; // @[LZD.scala 39:14]
  wire  _T_41; // @[LZD.scala 39:21]
  wire  _T_42; // @[LZD.scala 39:30]
  wire  _T_43; // @[LZD.scala 39:27]
  wire  _T_44; // @[LZD.scala 39:25]
  wire [1:0] _T_45; // @[Cat.scala 29:58]
  wire [1:0] _T_46; // @[LZD.scala 44:32]
  wire  _T_47; // @[LZD.scala 39:14]
  wire  _T_48; // @[LZD.scala 39:21]
  wire  _T_49; // @[LZD.scala 39:30]
  wire  _T_50; // @[LZD.scala 39:27]
  wire  _T_51; // @[LZD.scala 39:25]
  wire [1:0] _T_52; // @[Cat.scala 29:58]
  wire  _T_53; // @[Shift.scala 12:21]
  wire  _T_54; // @[Shift.scala 12:21]
  wire  _T_55; // @[LZD.scala 49:16]
  wire  _T_56; // @[LZD.scala 49:27]
  wire  _T_57; // @[LZD.scala 49:25]
  wire  _T_58; // @[LZD.scala 49:47]
  wire  _T_59; // @[LZD.scala 49:59]
  wire  _T_60; // @[LZD.scala 49:35]
  wire [2:0] _T_62; // @[Cat.scala 29:58]
  wire  _T_63; // @[Shift.scala 12:21]
  wire  _T_64; // @[Shift.scala 12:21]
  wire  _T_65; // @[LZD.scala 49:16]
  wire  _T_66; // @[LZD.scala 49:27]
  wire  _T_67; // @[LZD.scala 49:25]
  wire [1:0] _T_68; // @[LZD.scala 49:47]
  wire [1:0] _T_69; // @[LZD.scala 49:59]
  wire [1:0] _T_70; // @[LZD.scala 49:35]
  wire [3:0] _T_72; // @[Cat.scala 29:58]
  wire [7:0] _T_73; // @[LZD.scala 44:32]
  wire [3:0] _T_74; // @[LZD.scala 43:32]
  wire [1:0] _T_75; // @[LZD.scala 43:32]
  wire  _T_76; // @[LZD.scala 39:14]
  wire  _T_77; // @[LZD.scala 39:21]
  wire  _T_78; // @[LZD.scala 39:30]
  wire  _T_79; // @[LZD.scala 39:27]
  wire  _T_80; // @[LZD.scala 39:25]
  wire [1:0] _T_81; // @[Cat.scala 29:58]
  wire [1:0] _T_82; // @[LZD.scala 44:32]
  wire  _T_83; // @[LZD.scala 39:14]
  wire  _T_84; // @[LZD.scala 39:21]
  wire  _T_85; // @[LZD.scala 39:30]
  wire  _T_86; // @[LZD.scala 39:27]
  wire  _T_87; // @[LZD.scala 39:25]
  wire [1:0] _T_88; // @[Cat.scala 29:58]
  wire  _T_89; // @[Shift.scala 12:21]
  wire  _T_90; // @[Shift.scala 12:21]
  wire  _T_91; // @[LZD.scala 49:16]
  wire  _T_92; // @[LZD.scala 49:27]
  wire  _T_93; // @[LZD.scala 49:25]
  wire  _T_94; // @[LZD.scala 49:47]
  wire  _T_95; // @[LZD.scala 49:59]
  wire  _T_96; // @[LZD.scala 49:35]
  wire [2:0] _T_98; // @[Cat.scala 29:58]
  wire [3:0] _T_99; // @[LZD.scala 44:32]
  wire [1:0] _T_100; // @[LZD.scala 43:32]
  wire  _T_101; // @[LZD.scala 39:14]
  wire  _T_102; // @[LZD.scala 39:21]
  wire  _T_103; // @[LZD.scala 39:30]
  wire  _T_104; // @[LZD.scala 39:27]
  wire  _T_105; // @[LZD.scala 39:25]
  wire [1:0] _T_106; // @[Cat.scala 29:58]
  wire [1:0] _T_107; // @[LZD.scala 44:32]
  wire  _T_108; // @[LZD.scala 39:14]
  wire  _T_109; // @[LZD.scala 39:21]
  wire  _T_110; // @[LZD.scala 39:30]
  wire  _T_111; // @[LZD.scala 39:27]
  wire  _T_112; // @[LZD.scala 39:25]
  wire [1:0] _T_113; // @[Cat.scala 29:58]
  wire  _T_114; // @[Shift.scala 12:21]
  wire  _T_115; // @[Shift.scala 12:21]
  wire  _T_116; // @[LZD.scala 49:16]
  wire  _T_117; // @[LZD.scala 49:27]
  wire  _T_118; // @[LZD.scala 49:25]
  wire  _T_119; // @[LZD.scala 49:47]
  wire  _T_120; // @[LZD.scala 49:59]
  wire  _T_121; // @[LZD.scala 49:35]
  wire [2:0] _T_123; // @[Cat.scala 29:58]
  wire  _T_124; // @[Shift.scala 12:21]
  wire  _T_125; // @[Shift.scala 12:21]
  wire  _T_126; // @[LZD.scala 49:16]
  wire  _T_127; // @[LZD.scala 49:27]
  wire  _T_128; // @[LZD.scala 49:25]
  wire [1:0] _T_129; // @[LZD.scala 49:47]
  wire [1:0] _T_130; // @[LZD.scala 49:59]
  wire [1:0] _T_131; // @[LZD.scala 49:35]
  wire [3:0] _T_133; // @[Cat.scala 29:58]
  wire  _T_134; // @[Shift.scala 12:21]
  wire  _T_135; // @[Shift.scala 12:21]
  wire  _T_136; // @[LZD.scala 49:16]
  wire  _T_137; // @[LZD.scala 49:27]
  wire  _T_138; // @[LZD.scala 49:25]
  wire [2:0] _T_139; // @[LZD.scala 49:47]
  wire [2:0] _T_140; // @[LZD.scala 49:59]
  wire [2:0] _T_141; // @[LZD.scala 49:35]
  wire [4:0] _T_143; // @[Cat.scala 29:58]
  wire [15:0] _T_144; // @[LZD.scala 44:32]
  wire [7:0] _T_145; // @[LZD.scala 43:32]
  wire [3:0] _T_146; // @[LZD.scala 43:32]
  wire [1:0] _T_147; // @[LZD.scala 43:32]
  wire  _T_148; // @[LZD.scala 39:14]
  wire  _T_149; // @[LZD.scala 39:21]
  wire  _T_150; // @[LZD.scala 39:30]
  wire  _T_151; // @[LZD.scala 39:27]
  wire  _T_152; // @[LZD.scala 39:25]
  wire [1:0] _T_153; // @[Cat.scala 29:58]
  wire [1:0] _T_154; // @[LZD.scala 44:32]
  wire  _T_155; // @[LZD.scala 39:14]
  wire  _T_156; // @[LZD.scala 39:21]
  wire  _T_157; // @[LZD.scala 39:30]
  wire  _T_158; // @[LZD.scala 39:27]
  wire  _T_159; // @[LZD.scala 39:25]
  wire [1:0] _T_160; // @[Cat.scala 29:58]
  wire  _T_161; // @[Shift.scala 12:21]
  wire  _T_162; // @[Shift.scala 12:21]
  wire  _T_163; // @[LZD.scala 49:16]
  wire  _T_164; // @[LZD.scala 49:27]
  wire  _T_165; // @[LZD.scala 49:25]
  wire  _T_166; // @[LZD.scala 49:47]
  wire  _T_167; // @[LZD.scala 49:59]
  wire  _T_168; // @[LZD.scala 49:35]
  wire [2:0] _T_170; // @[Cat.scala 29:58]
  wire [3:0] _T_171; // @[LZD.scala 44:32]
  wire [1:0] _T_172; // @[LZD.scala 43:32]
  wire  _T_173; // @[LZD.scala 39:14]
  wire  _T_174; // @[LZD.scala 39:21]
  wire  _T_175; // @[LZD.scala 39:30]
  wire  _T_176; // @[LZD.scala 39:27]
  wire  _T_177; // @[LZD.scala 39:25]
  wire [1:0] _T_178; // @[Cat.scala 29:58]
  wire [1:0] _T_179; // @[LZD.scala 44:32]
  wire  _T_180; // @[LZD.scala 39:14]
  wire  _T_181; // @[LZD.scala 39:21]
  wire  _T_182; // @[LZD.scala 39:30]
  wire  _T_183; // @[LZD.scala 39:27]
  wire  _T_184; // @[LZD.scala 39:25]
  wire [1:0] _T_185; // @[Cat.scala 29:58]
  wire  _T_186; // @[Shift.scala 12:21]
  wire  _T_187; // @[Shift.scala 12:21]
  wire  _T_188; // @[LZD.scala 49:16]
  wire  _T_189; // @[LZD.scala 49:27]
  wire  _T_190; // @[LZD.scala 49:25]
  wire  _T_191; // @[LZD.scala 49:47]
  wire  _T_192; // @[LZD.scala 49:59]
  wire  _T_193; // @[LZD.scala 49:35]
  wire [2:0] _T_195; // @[Cat.scala 29:58]
  wire  _T_196; // @[Shift.scala 12:21]
  wire  _T_197; // @[Shift.scala 12:21]
  wire  _T_198; // @[LZD.scala 49:16]
  wire  _T_199; // @[LZD.scala 49:27]
  wire  _T_200; // @[LZD.scala 49:25]
  wire [1:0] _T_201; // @[LZD.scala 49:47]
  wire [1:0] _T_202; // @[LZD.scala 49:59]
  wire [1:0] _T_203; // @[LZD.scala 49:35]
  wire [3:0] _T_205; // @[Cat.scala 29:58]
  wire [7:0] _T_206; // @[LZD.scala 44:32]
  wire [3:0] _T_207; // @[LZD.scala 43:32]
  wire [1:0] _T_208; // @[LZD.scala 43:32]
  wire  _T_209; // @[LZD.scala 39:14]
  wire  _T_210; // @[LZD.scala 39:21]
  wire  _T_211; // @[LZD.scala 39:30]
  wire  _T_212; // @[LZD.scala 39:27]
  wire  _T_213; // @[LZD.scala 39:25]
  wire [1:0] _T_214; // @[Cat.scala 29:58]
  wire [1:0] _T_215; // @[LZD.scala 44:32]
  wire  _T_216; // @[LZD.scala 39:14]
  wire  _T_217; // @[LZD.scala 39:21]
  wire  _T_218; // @[LZD.scala 39:30]
  wire  _T_219; // @[LZD.scala 39:27]
  wire  _T_220; // @[LZD.scala 39:25]
  wire [1:0] _T_221; // @[Cat.scala 29:58]
  wire  _T_222; // @[Shift.scala 12:21]
  wire  _T_223; // @[Shift.scala 12:21]
  wire  _T_224; // @[LZD.scala 49:16]
  wire  _T_225; // @[LZD.scala 49:27]
  wire  _T_226; // @[LZD.scala 49:25]
  wire  _T_227; // @[LZD.scala 49:47]
  wire  _T_228; // @[LZD.scala 49:59]
  wire  _T_229; // @[LZD.scala 49:35]
  wire [2:0] _T_231; // @[Cat.scala 29:58]
  wire [3:0] _T_232; // @[LZD.scala 44:32]
  wire [1:0] _T_233; // @[LZD.scala 43:32]
  wire  _T_234; // @[LZD.scala 39:14]
  wire  _T_235; // @[LZD.scala 39:21]
  wire  _T_236; // @[LZD.scala 39:30]
  wire  _T_237; // @[LZD.scala 39:27]
  wire  _T_238; // @[LZD.scala 39:25]
  wire [1:0] _T_239; // @[Cat.scala 29:58]
  wire [1:0] _T_240; // @[LZD.scala 44:32]
  wire  _T_241; // @[LZD.scala 39:14]
  wire  _T_242; // @[LZD.scala 39:21]
  wire  _T_243; // @[LZD.scala 39:30]
  wire  _T_244; // @[LZD.scala 39:27]
  wire  _T_245; // @[LZD.scala 39:25]
  wire [1:0] _T_246; // @[Cat.scala 29:58]
  wire  _T_247; // @[Shift.scala 12:21]
  wire  _T_248; // @[Shift.scala 12:21]
  wire  _T_249; // @[LZD.scala 49:16]
  wire  _T_250; // @[LZD.scala 49:27]
  wire  _T_251; // @[LZD.scala 49:25]
  wire  _T_252; // @[LZD.scala 49:47]
  wire  _T_253; // @[LZD.scala 49:59]
  wire  _T_254; // @[LZD.scala 49:35]
  wire [2:0] _T_256; // @[Cat.scala 29:58]
  wire  _T_257; // @[Shift.scala 12:21]
  wire  _T_258; // @[Shift.scala 12:21]
  wire  _T_259; // @[LZD.scala 49:16]
  wire  _T_260; // @[LZD.scala 49:27]
  wire  _T_261; // @[LZD.scala 49:25]
  wire [1:0] _T_262; // @[LZD.scala 49:47]
  wire [1:0] _T_263; // @[LZD.scala 49:59]
  wire [1:0] _T_264; // @[LZD.scala 49:35]
  wire [3:0] _T_266; // @[Cat.scala 29:58]
  wire  _T_267; // @[Shift.scala 12:21]
  wire  _T_268; // @[Shift.scala 12:21]
  wire  _T_269; // @[LZD.scala 49:16]
  wire  _T_270; // @[LZD.scala 49:27]
  wire  _T_271; // @[LZD.scala 49:25]
  wire [2:0] _T_272; // @[LZD.scala 49:47]
  wire [2:0] _T_273; // @[LZD.scala 49:59]
  wire [2:0] _T_274; // @[LZD.scala 49:35]
  wire [4:0] _T_276; // @[Cat.scala 29:58]
  wire  _T_277; // @[Shift.scala 12:21]
  wire  _T_278; // @[Shift.scala 12:21]
  wire  _T_279; // @[LZD.scala 49:16]
  wire  _T_280; // @[LZD.scala 49:27]
  wire  _T_281; // @[LZD.scala 49:25]
  wire [3:0] _T_282; // @[LZD.scala 49:47]
  wire [3:0] _T_283; // @[LZD.scala 49:59]
  wire [3:0] _T_284; // @[LZD.scala 49:35]
  wire [5:0] _T_286; // @[Cat.scala 29:58]
  wire [30:0] _T_287; // @[LZD.scala 44:32]
  wire [15:0] _T_288; // @[LZD.scala 43:32]
  wire [7:0] _T_289; // @[LZD.scala 43:32]
  wire [3:0] _T_290; // @[LZD.scala 43:32]
  wire [1:0] _T_291; // @[LZD.scala 43:32]
  wire  _T_292; // @[LZD.scala 39:14]
  wire  _T_293; // @[LZD.scala 39:21]
  wire  _T_294; // @[LZD.scala 39:30]
  wire  _T_295; // @[LZD.scala 39:27]
  wire  _T_296; // @[LZD.scala 39:25]
  wire [1:0] _T_297; // @[Cat.scala 29:58]
  wire [1:0] _T_298; // @[LZD.scala 44:32]
  wire  _T_299; // @[LZD.scala 39:14]
  wire  _T_300; // @[LZD.scala 39:21]
  wire  _T_301; // @[LZD.scala 39:30]
  wire  _T_302; // @[LZD.scala 39:27]
  wire  _T_303; // @[LZD.scala 39:25]
  wire [1:0] _T_304; // @[Cat.scala 29:58]
  wire  _T_305; // @[Shift.scala 12:21]
  wire  _T_306; // @[Shift.scala 12:21]
  wire  _T_307; // @[LZD.scala 49:16]
  wire  _T_308; // @[LZD.scala 49:27]
  wire  _T_309; // @[LZD.scala 49:25]
  wire  _T_310; // @[LZD.scala 49:47]
  wire  _T_311; // @[LZD.scala 49:59]
  wire  _T_312; // @[LZD.scala 49:35]
  wire [2:0] _T_314; // @[Cat.scala 29:58]
  wire [3:0] _T_315; // @[LZD.scala 44:32]
  wire [1:0] _T_316; // @[LZD.scala 43:32]
  wire  _T_317; // @[LZD.scala 39:14]
  wire  _T_318; // @[LZD.scala 39:21]
  wire  _T_319; // @[LZD.scala 39:30]
  wire  _T_320; // @[LZD.scala 39:27]
  wire  _T_321; // @[LZD.scala 39:25]
  wire [1:0] _T_322; // @[Cat.scala 29:58]
  wire [1:0] _T_323; // @[LZD.scala 44:32]
  wire  _T_324; // @[LZD.scala 39:14]
  wire  _T_325; // @[LZD.scala 39:21]
  wire  _T_326; // @[LZD.scala 39:30]
  wire  _T_327; // @[LZD.scala 39:27]
  wire  _T_328; // @[LZD.scala 39:25]
  wire [1:0] _T_329; // @[Cat.scala 29:58]
  wire  _T_330; // @[Shift.scala 12:21]
  wire  _T_331; // @[Shift.scala 12:21]
  wire  _T_332; // @[LZD.scala 49:16]
  wire  _T_333; // @[LZD.scala 49:27]
  wire  _T_334; // @[LZD.scala 49:25]
  wire  _T_335; // @[LZD.scala 49:47]
  wire  _T_336; // @[LZD.scala 49:59]
  wire  _T_337; // @[LZD.scala 49:35]
  wire [2:0] _T_339; // @[Cat.scala 29:58]
  wire  _T_340; // @[Shift.scala 12:21]
  wire  _T_341; // @[Shift.scala 12:21]
  wire  _T_342; // @[LZD.scala 49:16]
  wire  _T_343; // @[LZD.scala 49:27]
  wire  _T_344; // @[LZD.scala 49:25]
  wire [1:0] _T_345; // @[LZD.scala 49:47]
  wire [1:0] _T_346; // @[LZD.scala 49:59]
  wire [1:0] _T_347; // @[LZD.scala 49:35]
  wire [3:0] _T_349; // @[Cat.scala 29:58]
  wire [7:0] _T_350; // @[LZD.scala 44:32]
  wire [3:0] _T_351; // @[LZD.scala 43:32]
  wire [1:0] _T_352; // @[LZD.scala 43:32]
  wire  _T_353; // @[LZD.scala 39:14]
  wire  _T_354; // @[LZD.scala 39:21]
  wire  _T_355; // @[LZD.scala 39:30]
  wire  _T_356; // @[LZD.scala 39:27]
  wire  _T_357; // @[LZD.scala 39:25]
  wire [1:0] _T_358; // @[Cat.scala 29:58]
  wire [1:0] _T_359; // @[LZD.scala 44:32]
  wire  _T_360; // @[LZD.scala 39:14]
  wire  _T_361; // @[LZD.scala 39:21]
  wire  _T_362; // @[LZD.scala 39:30]
  wire  _T_363; // @[LZD.scala 39:27]
  wire  _T_364; // @[LZD.scala 39:25]
  wire [1:0] _T_365; // @[Cat.scala 29:58]
  wire  _T_366; // @[Shift.scala 12:21]
  wire  _T_367; // @[Shift.scala 12:21]
  wire  _T_368; // @[LZD.scala 49:16]
  wire  _T_369; // @[LZD.scala 49:27]
  wire  _T_370; // @[LZD.scala 49:25]
  wire  _T_371; // @[LZD.scala 49:47]
  wire  _T_372; // @[LZD.scala 49:59]
  wire  _T_373; // @[LZD.scala 49:35]
  wire [2:0] _T_375; // @[Cat.scala 29:58]
  wire [3:0] _T_376; // @[LZD.scala 44:32]
  wire [1:0] _T_377; // @[LZD.scala 43:32]
  wire  _T_378; // @[LZD.scala 39:14]
  wire  _T_379; // @[LZD.scala 39:21]
  wire  _T_380; // @[LZD.scala 39:30]
  wire  _T_381; // @[LZD.scala 39:27]
  wire  _T_382; // @[LZD.scala 39:25]
  wire [1:0] _T_383; // @[Cat.scala 29:58]
  wire [1:0] _T_384; // @[LZD.scala 44:32]
  wire  _T_385; // @[LZD.scala 39:14]
  wire  _T_386; // @[LZD.scala 39:21]
  wire  _T_387; // @[LZD.scala 39:30]
  wire  _T_388; // @[LZD.scala 39:27]
  wire  _T_389; // @[LZD.scala 39:25]
  wire [1:0] _T_390; // @[Cat.scala 29:58]
  wire  _T_391; // @[Shift.scala 12:21]
  wire  _T_392; // @[Shift.scala 12:21]
  wire  _T_393; // @[LZD.scala 49:16]
  wire  _T_394; // @[LZD.scala 49:27]
  wire  _T_395; // @[LZD.scala 49:25]
  wire  _T_396; // @[LZD.scala 49:47]
  wire  _T_397; // @[LZD.scala 49:59]
  wire  _T_398; // @[LZD.scala 49:35]
  wire [2:0] _T_400; // @[Cat.scala 29:58]
  wire  _T_401; // @[Shift.scala 12:21]
  wire  _T_402; // @[Shift.scala 12:21]
  wire  _T_403; // @[LZD.scala 49:16]
  wire  _T_404; // @[LZD.scala 49:27]
  wire  _T_405; // @[LZD.scala 49:25]
  wire [1:0] _T_406; // @[LZD.scala 49:47]
  wire [1:0] _T_407; // @[LZD.scala 49:59]
  wire [1:0] _T_408; // @[LZD.scala 49:35]
  wire [3:0] _T_410; // @[Cat.scala 29:58]
  wire  _T_411; // @[Shift.scala 12:21]
  wire  _T_412; // @[Shift.scala 12:21]
  wire  _T_413; // @[LZD.scala 49:16]
  wire  _T_414; // @[LZD.scala 49:27]
  wire  _T_415; // @[LZD.scala 49:25]
  wire [2:0] _T_416; // @[LZD.scala 49:47]
  wire [2:0] _T_417; // @[LZD.scala 49:59]
  wire [2:0] _T_418; // @[LZD.scala 49:35]
  wire [4:0] _T_420; // @[Cat.scala 29:58]
  wire [14:0] _T_421; // @[LZD.scala 44:32]
  wire [7:0] _T_422; // @[LZD.scala 43:32]
  wire [3:0] _T_423; // @[LZD.scala 43:32]
  wire [1:0] _T_424; // @[LZD.scala 43:32]
  wire  _T_425; // @[LZD.scala 39:14]
  wire  _T_426; // @[LZD.scala 39:21]
  wire  _T_427; // @[LZD.scala 39:30]
  wire  _T_428; // @[LZD.scala 39:27]
  wire  _T_429; // @[LZD.scala 39:25]
  wire [1:0] _T_430; // @[Cat.scala 29:58]
  wire [1:0] _T_431; // @[LZD.scala 44:32]
  wire  _T_432; // @[LZD.scala 39:14]
  wire  _T_433; // @[LZD.scala 39:21]
  wire  _T_434; // @[LZD.scala 39:30]
  wire  _T_435; // @[LZD.scala 39:27]
  wire  _T_436; // @[LZD.scala 39:25]
  wire [1:0] _T_437; // @[Cat.scala 29:58]
  wire  _T_438; // @[Shift.scala 12:21]
  wire  _T_439; // @[Shift.scala 12:21]
  wire  _T_440; // @[LZD.scala 49:16]
  wire  _T_441; // @[LZD.scala 49:27]
  wire  _T_442; // @[LZD.scala 49:25]
  wire  _T_443; // @[LZD.scala 49:47]
  wire  _T_444; // @[LZD.scala 49:59]
  wire  _T_445; // @[LZD.scala 49:35]
  wire [2:0] _T_447; // @[Cat.scala 29:58]
  wire [3:0] _T_448; // @[LZD.scala 44:32]
  wire [1:0] _T_449; // @[LZD.scala 43:32]
  wire  _T_450; // @[LZD.scala 39:14]
  wire  _T_451; // @[LZD.scala 39:21]
  wire  _T_452; // @[LZD.scala 39:30]
  wire  _T_453; // @[LZD.scala 39:27]
  wire  _T_454; // @[LZD.scala 39:25]
  wire [1:0] _T_455; // @[Cat.scala 29:58]
  wire [1:0] _T_456; // @[LZD.scala 44:32]
  wire  _T_457; // @[LZD.scala 39:14]
  wire  _T_458; // @[LZD.scala 39:21]
  wire  _T_459; // @[LZD.scala 39:30]
  wire  _T_460; // @[LZD.scala 39:27]
  wire  _T_461; // @[LZD.scala 39:25]
  wire [1:0] _T_462; // @[Cat.scala 29:58]
  wire  _T_463; // @[Shift.scala 12:21]
  wire  _T_464; // @[Shift.scala 12:21]
  wire  _T_465; // @[LZD.scala 49:16]
  wire  _T_466; // @[LZD.scala 49:27]
  wire  _T_467; // @[LZD.scala 49:25]
  wire  _T_468; // @[LZD.scala 49:47]
  wire  _T_469; // @[LZD.scala 49:59]
  wire  _T_470; // @[LZD.scala 49:35]
  wire [2:0] _T_472; // @[Cat.scala 29:58]
  wire  _T_473; // @[Shift.scala 12:21]
  wire  _T_474; // @[Shift.scala 12:21]
  wire  _T_475; // @[LZD.scala 49:16]
  wire  _T_476; // @[LZD.scala 49:27]
  wire  _T_477; // @[LZD.scala 49:25]
  wire [1:0] _T_478; // @[LZD.scala 49:47]
  wire [1:0] _T_479; // @[LZD.scala 49:59]
  wire [1:0] _T_480; // @[LZD.scala 49:35]
  wire [3:0] _T_482; // @[Cat.scala 29:58]
  wire [6:0] _T_483; // @[LZD.scala 44:32]
  wire [3:0] _T_484; // @[LZD.scala 43:32]
  wire [1:0] _T_485; // @[LZD.scala 43:32]
  wire  _T_486; // @[LZD.scala 39:14]
  wire  _T_487; // @[LZD.scala 39:21]
  wire  _T_488; // @[LZD.scala 39:30]
  wire  _T_489; // @[LZD.scala 39:27]
  wire  _T_490; // @[LZD.scala 39:25]
  wire [1:0] _T_491; // @[Cat.scala 29:58]
  wire [1:0] _T_492; // @[LZD.scala 44:32]
  wire  _T_493; // @[LZD.scala 39:14]
  wire  _T_494; // @[LZD.scala 39:21]
  wire  _T_495; // @[LZD.scala 39:30]
  wire  _T_496; // @[LZD.scala 39:27]
  wire  _T_497; // @[LZD.scala 39:25]
  wire [1:0] _T_498; // @[Cat.scala 29:58]
  wire  _T_499; // @[Shift.scala 12:21]
  wire  _T_500; // @[Shift.scala 12:21]
  wire  _T_501; // @[LZD.scala 49:16]
  wire  _T_502; // @[LZD.scala 49:27]
  wire  _T_503; // @[LZD.scala 49:25]
  wire  _T_504; // @[LZD.scala 49:47]
  wire  _T_505; // @[LZD.scala 49:59]
  wire  _T_506; // @[LZD.scala 49:35]
  wire [2:0] _T_508; // @[Cat.scala 29:58]
  wire [2:0] _T_509; // @[LZD.scala 44:32]
  wire [1:0] _T_510; // @[LZD.scala 43:32]
  wire  _T_511; // @[LZD.scala 39:14]
  wire  _T_512; // @[LZD.scala 39:21]
  wire  _T_513; // @[LZD.scala 39:30]
  wire  _T_514; // @[LZD.scala 39:27]
  wire  _T_515; // @[LZD.scala 39:25]
  wire [1:0] _T_516; // @[Cat.scala 29:58]
  wire  _T_517; // @[LZD.scala 44:32]
  wire  _T_519; // @[Shift.scala 12:21]
  wire  _T_521; // @[LZD.scala 55:32]
  wire  _T_522; // @[LZD.scala 55:20]
  wire [1:0] _T_523; // @[Cat.scala 29:58]
  wire  _T_524; // @[Shift.scala 12:21]
  wire [1:0] _T_526; // @[LZD.scala 55:32]
  wire [1:0] _T_527; // @[LZD.scala 55:20]
  wire [2:0] _T_528; // @[Cat.scala 29:58]
  wire  _T_529; // @[Shift.scala 12:21]
  wire [2:0] _T_531; // @[LZD.scala 55:32]
  wire [2:0] _T_532; // @[LZD.scala 55:20]
  wire [3:0] _T_533; // @[Cat.scala 29:58]
  wire  _T_534; // @[Shift.scala 12:21]
  wire [3:0] _T_536; // @[LZD.scala 55:32]
  wire [3:0] _T_537; // @[LZD.scala 55:20]
  wire [4:0] _T_538; // @[Cat.scala 29:58]
  wire  _T_539; // @[Shift.scala 12:21]
  wire [4:0] _T_541; // @[LZD.scala 55:32]
  wire [4:0] _T_542; // @[LZD.scala 55:20]
  wire [6:0] scaleBias; // @[Cat.scala 29:58]
  wire [6:0] _T_543; // @[QuireToPosit.scala 61:53]
  wire [7:0] _GEN_2; // @[QuireToPosit.scala 61:41]
  wire [7:0] _T_545; // @[QuireToPosit.scala 61:41]
  wire [7:0] realScale; // @[QuireToPosit.scala 61:41]
  wire  underflow; // @[QuireToPosit.scala 62:41]
  wire  overflow; // @[QuireToPosit.scala 63:35]
  wire [7:0] _T_546; // @[Mux.scala 87:16]
  wire [7:0] _T_547; // @[Mux.scala 87:16]
  wire  _T_548; // @[Abs.scala 10:21]
  wire [7:0] _T_550; // @[Bitwise.scala 71:12]
  wire [7:0] _T_551; // @[Abs.scala 10:31]
  wire [7:0] _T_552; // @[Abs.scala 10:26]
  wire [7:0] _GEN_3; // @[Abs.scala 10:39]
  wire [7:0] absRealScale; // @[Abs.scala 10:39]
  wire  _T_555; // @[Shift.scala 16:24]
  wire [5:0] _T_556; // @[Shift.scala 17:37]
  wire  _T_557; // @[Shift.scala 12:21]
  wire [31:0] _T_558; // @[Shift.scala 64:52]
  wire [63:0] _T_560; // @[Cat.scala 29:58]
  wire [63:0] _T_561; // @[Shift.scala 64:27]
  wire [4:0] _T_562; // @[Shift.scala 66:70]
  wire  _T_563; // @[Shift.scala 12:21]
  wire [47:0] _T_564; // @[Shift.scala 64:52]
  wire [63:0] _T_566; // @[Cat.scala 29:58]
  wire [63:0] _T_567; // @[Shift.scala 64:27]
  wire [3:0] _T_568; // @[Shift.scala 66:70]
  wire  _T_569; // @[Shift.scala 12:21]
  wire [55:0] _T_570; // @[Shift.scala 64:52]
  wire [63:0] _T_572; // @[Cat.scala 29:58]
  wire [63:0] _T_573; // @[Shift.scala 64:27]
  wire [2:0] _T_574; // @[Shift.scala 66:70]
  wire  _T_575; // @[Shift.scala 12:21]
  wire [59:0] _T_576; // @[Shift.scala 64:52]
  wire [63:0] _T_578; // @[Cat.scala 29:58]
  wire [63:0] _T_579; // @[Shift.scala 64:27]
  wire [1:0] _T_580; // @[Shift.scala 66:70]
  wire  _T_581; // @[Shift.scala 12:21]
  wire [61:0] _T_582; // @[Shift.scala 64:52]
  wire [63:0] _T_584; // @[Cat.scala 29:58]
  wire [63:0] _T_585; // @[Shift.scala 64:27]
  wire  _T_586; // @[Shift.scala 66:70]
  wire [62:0] _T_588; // @[Shift.scala 64:52]
  wire [63:0] _T_589; // @[Cat.scala 29:58]
  wire [63:0] _T_590; // @[Shift.scala 64:27]
  wire [63:0] quireLeftShift; // @[Shift.scala 16:10]
  wire [31:0] _T_595; // @[Shift.scala 77:66]
  wire [63:0] _T_596; // @[Cat.scala 29:58]
  wire [63:0] _T_597; // @[Shift.scala 77:22]
  wire [47:0] _T_601; // @[Shift.scala 77:66]
  wire [63:0] _T_602; // @[Cat.scala 29:58]
  wire [63:0] _T_603; // @[Shift.scala 77:22]
  wire [55:0] _T_607; // @[Shift.scala 77:66]
  wire [63:0] _T_608; // @[Cat.scala 29:58]
  wire [63:0] _T_609; // @[Shift.scala 77:22]
  wire [59:0] _T_613; // @[Shift.scala 77:66]
  wire [63:0] _T_614; // @[Cat.scala 29:58]
  wire [63:0] _T_615; // @[Shift.scala 77:22]
  wire [61:0] _T_619; // @[Shift.scala 77:66]
  wire [63:0] _T_620; // @[Cat.scala 29:58]
  wire [63:0] _T_621; // @[Shift.scala 77:22]
  wire [62:0] _T_624; // @[Shift.scala 77:66]
  wire [63:0] _T_625; // @[Cat.scala 29:58]
  wire [63:0] _T_626; // @[Shift.scala 77:22]
  wire [63:0] quireRightShift; // @[Shift.scala 27:10]
  wire [5:0] _T_628; // @[QuireToPosit.scala 89:49]
  wire [17:0] _T_629; // @[QuireToPosit.scala 90:127]
  wire  _T_630; // @[QuireToPosit.scala 90:154]
  wire [6:0] realFGRSTmp1; // @[Cat.scala 29:58]
  wire [5:0] _T_631; // @[QuireToPosit.scala 91:50]
  wire [17:0] _T_632; // @[QuireToPosit.scala 92:128]
  wire  _T_633; // @[QuireToPosit.scala 92:155]
  wire [6:0] realFGRSTmp2; // @[Cat.scala 29:58]
  wire [6:0] realFGRS; // @[QuireToPosit.scala 93:34]
  wire [3:0] outRawFloat_fraction; // @[QuireToPosit.scala 95:46]
  wire [2:0] outRawFloat_grs; // @[QuireToPosit.scala 96:46]
  wire [4:0] _GEN_4; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  wire [4:0] outRawFloat_scale; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  wire  _T_638; // @[convert.scala 46:61]
  wire  _T_639; // @[convert.scala 46:52]
  wire  _T_641; // @[convert.scala 46:42]
  wire [3:0] _T_642; // @[convert.scala 48:34]
  wire  _T_643; // @[convert.scala 49:36]
  wire [3:0] _T_645; // @[convert.scala 50:36]
  wire [3:0] _T_646; // @[convert.scala 50:36]
  wire [3:0] _T_647; // @[convert.scala 50:28]
  wire  _T_648; // @[convert.scala 51:31]
  wire  _T_649; // @[convert.scala 52:43]
  wire [9:0] _T_653; // @[Cat.scala 29:58]
  wire [3:0] _T_654; // @[Shift.scala 39:17]
  wire  _T_655; // @[Shift.scala 39:24]
  wire [1:0] _T_657; // @[Shift.scala 90:30]
  wire [7:0] _T_658; // @[Shift.scala 90:48]
  wire  _T_659; // @[Shift.scala 90:57]
  wire [1:0] _GEN_5; // @[Shift.scala 90:39]
  wire [1:0] _T_660; // @[Shift.scala 90:39]
  wire  _T_661; // @[Shift.scala 12:21]
  wire  _T_662; // @[Shift.scala 12:21]
  wire [7:0] _T_664; // @[Bitwise.scala 71:12]
  wire [9:0] _T_665; // @[Cat.scala 29:58]
  wire [9:0] _T_666; // @[Shift.scala 91:22]
  wire [2:0] _T_667; // @[Shift.scala 92:77]
  wire [5:0] _T_668; // @[Shift.scala 90:30]
  wire [3:0] _T_669; // @[Shift.scala 90:48]
  wire  _T_670; // @[Shift.scala 90:57]
  wire [5:0] _GEN_6; // @[Shift.scala 90:39]
  wire [5:0] _T_671; // @[Shift.scala 90:39]
  wire  _T_672; // @[Shift.scala 12:21]
  wire  _T_673; // @[Shift.scala 12:21]
  wire [3:0] _T_675; // @[Bitwise.scala 71:12]
  wire [9:0] _T_676; // @[Cat.scala 29:58]
  wire [9:0] _T_677; // @[Shift.scala 91:22]
  wire [1:0] _T_678; // @[Shift.scala 92:77]
  wire [7:0] _T_679; // @[Shift.scala 90:30]
  wire [1:0] _T_680; // @[Shift.scala 90:48]
  wire  _T_681; // @[Shift.scala 90:57]
  wire [7:0] _GEN_7; // @[Shift.scala 90:39]
  wire [7:0] _T_682; // @[Shift.scala 90:39]
  wire  _T_683; // @[Shift.scala 12:21]
  wire  _T_684; // @[Shift.scala 12:21]
  wire [1:0] _T_686; // @[Bitwise.scala 71:12]
  wire [9:0] _T_687; // @[Cat.scala 29:58]
  wire [9:0] _T_688; // @[Shift.scala 91:22]
  wire  _T_689; // @[Shift.scala 92:77]
  wire [8:0] _T_690; // @[Shift.scala 90:30]
  wire  _T_691; // @[Shift.scala 90:48]
  wire [8:0] _GEN_8; // @[Shift.scala 90:39]
  wire [8:0] _T_693; // @[Shift.scala 90:39]
  wire  _T_695; // @[Shift.scala 12:21]
  wire [9:0] _T_696; // @[Cat.scala 29:58]
  wire [9:0] _T_697; // @[Shift.scala 91:22]
  wire [9:0] _T_700; // @[Bitwise.scala 71:12]
  wire [9:0] _T_701; // @[Shift.scala 39:10]
  wire  _T_702; // @[convert.scala 55:31]
  wire  _T_703; // @[convert.scala 56:31]
  wire  _T_704; // @[convert.scala 57:31]
  wire  _T_705; // @[convert.scala 58:31]
  wire [6:0] _T_706; // @[convert.scala 59:69]
  wire  _T_707; // @[convert.scala 59:81]
  wire  _T_708; // @[convert.scala 59:50]
  wire  _T_710; // @[convert.scala 60:81]
  wire  _T_711; // @[convert.scala 61:44]
  wire  _T_712; // @[convert.scala 61:52]
  wire  _T_713; // @[convert.scala 61:36]
  wire  _T_714; // @[convert.scala 62:63]
  wire  _T_715; // @[convert.scala 62:103]
  wire  _T_716; // @[convert.scala 62:60]
  wire [6:0] _GEN_9; // @[convert.scala 63:56]
  wire [6:0] _T_719; // @[convert.scala 63:56]
  wire [7:0] _T_720; // @[Cat.scala 29:58]
  reg  _T_724; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [7:0] _T_728; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  assign _T = io_quireIn[62:0]; // @[QuireToPosit.scala 47:43]
  assign _T_1 = _T != 63'h0; // @[QuireToPosit.scala 47:47]
  assign tailIsZero = ~ _T_1; // @[QuireToPosit.scala 47:27]
  assign _T_2 = io_quireIn[63:63]; // @[QuireToPosit.scala 49:45]
  assign outRawFloat_isNaR = _T_2 & tailIsZero; // @[QuireToPosit.scala 49:49]
  assign _T_5 = ~ _T_2; // @[QuireToPosit.scala 50:31]
  assign outRawFloat_isZero = _T_5 & tailIsZero; // @[QuireToPosit.scala 50:51]
  assign _T_8 = io_quireIn[63:1]; // @[QuireToPosit.scala 58:41]
  assign _T_9 = io_quireIn[62:0]; // @[QuireToPosit.scala 58:68]
  assign quireXOR = _T_8 ^ _T_9; // @[QuireToPosit.scala 58:56]
  assign _T_10 = quireXOR[62:31]; // @[LZD.scala 43:32]
  assign _T_11 = _T_10[31:16]; // @[LZD.scala 43:32]
  assign _T_12 = _T_11[15:8]; // @[LZD.scala 43:32]
  assign _T_13 = _T_12[7:4]; // @[LZD.scala 43:32]
  assign _T_14 = _T_13[3:2]; // @[LZD.scala 43:32]
  assign _T_15 = _T_14 != 2'h0; // @[LZD.scala 39:14]
  assign _T_16 = _T_14[1]; // @[LZD.scala 39:21]
  assign _T_17 = _T_14[0]; // @[LZD.scala 39:30]
  assign _T_18 = ~ _T_17; // @[LZD.scala 39:27]
  assign _T_19 = _T_16 | _T_18; // @[LZD.scala 39:25]
  assign _T_20 = {_T_15,_T_19}; // @[Cat.scala 29:58]
  assign _T_21 = _T_13[1:0]; // @[LZD.scala 44:32]
  assign _T_22 = _T_21 != 2'h0; // @[LZD.scala 39:14]
  assign _T_23 = _T_21[1]; // @[LZD.scala 39:21]
  assign _T_24 = _T_21[0]; // @[LZD.scala 39:30]
  assign _T_25 = ~ _T_24; // @[LZD.scala 39:27]
  assign _T_26 = _T_23 | _T_25; // @[LZD.scala 39:25]
  assign _T_27 = {_T_22,_T_26}; // @[Cat.scala 29:58]
  assign _T_28 = _T_20[1]; // @[Shift.scala 12:21]
  assign _T_29 = _T_27[1]; // @[Shift.scala 12:21]
  assign _T_30 = _T_28 | _T_29; // @[LZD.scala 49:16]
  assign _T_31 = ~ _T_29; // @[LZD.scala 49:27]
  assign _T_32 = _T_28 | _T_31; // @[LZD.scala 49:25]
  assign _T_33 = _T_20[0:0]; // @[LZD.scala 49:47]
  assign _T_34 = _T_27[0:0]; // @[LZD.scala 49:59]
  assign _T_35 = _T_28 ? _T_33 : _T_34; // @[LZD.scala 49:35]
  assign _T_37 = {_T_30,_T_32,_T_35}; // @[Cat.scala 29:58]
  assign _T_38 = _T_12[3:0]; // @[LZD.scala 44:32]
  assign _T_39 = _T_38[3:2]; // @[LZD.scala 43:32]
  assign _T_40 = _T_39 != 2'h0; // @[LZD.scala 39:14]
  assign _T_41 = _T_39[1]; // @[LZD.scala 39:21]
  assign _T_42 = _T_39[0]; // @[LZD.scala 39:30]
  assign _T_43 = ~ _T_42; // @[LZD.scala 39:27]
  assign _T_44 = _T_41 | _T_43; // @[LZD.scala 39:25]
  assign _T_45 = {_T_40,_T_44}; // @[Cat.scala 29:58]
  assign _T_46 = _T_38[1:0]; // @[LZD.scala 44:32]
  assign _T_47 = _T_46 != 2'h0; // @[LZD.scala 39:14]
  assign _T_48 = _T_46[1]; // @[LZD.scala 39:21]
  assign _T_49 = _T_46[0]; // @[LZD.scala 39:30]
  assign _T_50 = ~ _T_49; // @[LZD.scala 39:27]
  assign _T_51 = _T_48 | _T_50; // @[LZD.scala 39:25]
  assign _T_52 = {_T_47,_T_51}; // @[Cat.scala 29:58]
  assign _T_53 = _T_45[1]; // @[Shift.scala 12:21]
  assign _T_54 = _T_52[1]; // @[Shift.scala 12:21]
  assign _T_55 = _T_53 | _T_54; // @[LZD.scala 49:16]
  assign _T_56 = ~ _T_54; // @[LZD.scala 49:27]
  assign _T_57 = _T_53 | _T_56; // @[LZD.scala 49:25]
  assign _T_58 = _T_45[0:0]; // @[LZD.scala 49:47]
  assign _T_59 = _T_52[0:0]; // @[LZD.scala 49:59]
  assign _T_60 = _T_53 ? _T_58 : _T_59; // @[LZD.scala 49:35]
  assign _T_62 = {_T_55,_T_57,_T_60}; // @[Cat.scala 29:58]
  assign _T_63 = _T_37[2]; // @[Shift.scala 12:21]
  assign _T_64 = _T_62[2]; // @[Shift.scala 12:21]
  assign _T_65 = _T_63 | _T_64; // @[LZD.scala 49:16]
  assign _T_66 = ~ _T_64; // @[LZD.scala 49:27]
  assign _T_67 = _T_63 | _T_66; // @[LZD.scala 49:25]
  assign _T_68 = _T_37[1:0]; // @[LZD.scala 49:47]
  assign _T_69 = _T_62[1:0]; // @[LZD.scala 49:59]
  assign _T_70 = _T_63 ? _T_68 : _T_69; // @[LZD.scala 49:35]
  assign _T_72 = {_T_65,_T_67,_T_70}; // @[Cat.scala 29:58]
  assign _T_73 = _T_11[7:0]; // @[LZD.scala 44:32]
  assign _T_74 = _T_73[7:4]; // @[LZD.scala 43:32]
  assign _T_75 = _T_74[3:2]; // @[LZD.scala 43:32]
  assign _T_76 = _T_75 != 2'h0; // @[LZD.scala 39:14]
  assign _T_77 = _T_75[1]; // @[LZD.scala 39:21]
  assign _T_78 = _T_75[0]; // @[LZD.scala 39:30]
  assign _T_79 = ~ _T_78; // @[LZD.scala 39:27]
  assign _T_80 = _T_77 | _T_79; // @[LZD.scala 39:25]
  assign _T_81 = {_T_76,_T_80}; // @[Cat.scala 29:58]
  assign _T_82 = _T_74[1:0]; // @[LZD.scala 44:32]
  assign _T_83 = _T_82 != 2'h0; // @[LZD.scala 39:14]
  assign _T_84 = _T_82[1]; // @[LZD.scala 39:21]
  assign _T_85 = _T_82[0]; // @[LZD.scala 39:30]
  assign _T_86 = ~ _T_85; // @[LZD.scala 39:27]
  assign _T_87 = _T_84 | _T_86; // @[LZD.scala 39:25]
  assign _T_88 = {_T_83,_T_87}; // @[Cat.scala 29:58]
  assign _T_89 = _T_81[1]; // @[Shift.scala 12:21]
  assign _T_90 = _T_88[1]; // @[Shift.scala 12:21]
  assign _T_91 = _T_89 | _T_90; // @[LZD.scala 49:16]
  assign _T_92 = ~ _T_90; // @[LZD.scala 49:27]
  assign _T_93 = _T_89 | _T_92; // @[LZD.scala 49:25]
  assign _T_94 = _T_81[0:0]; // @[LZD.scala 49:47]
  assign _T_95 = _T_88[0:0]; // @[LZD.scala 49:59]
  assign _T_96 = _T_89 ? _T_94 : _T_95; // @[LZD.scala 49:35]
  assign _T_98 = {_T_91,_T_93,_T_96}; // @[Cat.scala 29:58]
  assign _T_99 = _T_73[3:0]; // @[LZD.scala 44:32]
  assign _T_100 = _T_99[3:2]; // @[LZD.scala 43:32]
  assign _T_101 = _T_100 != 2'h0; // @[LZD.scala 39:14]
  assign _T_102 = _T_100[1]; // @[LZD.scala 39:21]
  assign _T_103 = _T_100[0]; // @[LZD.scala 39:30]
  assign _T_104 = ~ _T_103; // @[LZD.scala 39:27]
  assign _T_105 = _T_102 | _T_104; // @[LZD.scala 39:25]
  assign _T_106 = {_T_101,_T_105}; // @[Cat.scala 29:58]
  assign _T_107 = _T_99[1:0]; // @[LZD.scala 44:32]
  assign _T_108 = _T_107 != 2'h0; // @[LZD.scala 39:14]
  assign _T_109 = _T_107[1]; // @[LZD.scala 39:21]
  assign _T_110 = _T_107[0]; // @[LZD.scala 39:30]
  assign _T_111 = ~ _T_110; // @[LZD.scala 39:27]
  assign _T_112 = _T_109 | _T_111; // @[LZD.scala 39:25]
  assign _T_113 = {_T_108,_T_112}; // @[Cat.scala 29:58]
  assign _T_114 = _T_106[1]; // @[Shift.scala 12:21]
  assign _T_115 = _T_113[1]; // @[Shift.scala 12:21]
  assign _T_116 = _T_114 | _T_115; // @[LZD.scala 49:16]
  assign _T_117 = ~ _T_115; // @[LZD.scala 49:27]
  assign _T_118 = _T_114 | _T_117; // @[LZD.scala 49:25]
  assign _T_119 = _T_106[0:0]; // @[LZD.scala 49:47]
  assign _T_120 = _T_113[0:0]; // @[LZD.scala 49:59]
  assign _T_121 = _T_114 ? _T_119 : _T_120; // @[LZD.scala 49:35]
  assign _T_123 = {_T_116,_T_118,_T_121}; // @[Cat.scala 29:58]
  assign _T_124 = _T_98[2]; // @[Shift.scala 12:21]
  assign _T_125 = _T_123[2]; // @[Shift.scala 12:21]
  assign _T_126 = _T_124 | _T_125; // @[LZD.scala 49:16]
  assign _T_127 = ~ _T_125; // @[LZD.scala 49:27]
  assign _T_128 = _T_124 | _T_127; // @[LZD.scala 49:25]
  assign _T_129 = _T_98[1:0]; // @[LZD.scala 49:47]
  assign _T_130 = _T_123[1:0]; // @[LZD.scala 49:59]
  assign _T_131 = _T_124 ? _T_129 : _T_130; // @[LZD.scala 49:35]
  assign _T_133 = {_T_126,_T_128,_T_131}; // @[Cat.scala 29:58]
  assign _T_134 = _T_72[3]; // @[Shift.scala 12:21]
  assign _T_135 = _T_133[3]; // @[Shift.scala 12:21]
  assign _T_136 = _T_134 | _T_135; // @[LZD.scala 49:16]
  assign _T_137 = ~ _T_135; // @[LZD.scala 49:27]
  assign _T_138 = _T_134 | _T_137; // @[LZD.scala 49:25]
  assign _T_139 = _T_72[2:0]; // @[LZD.scala 49:47]
  assign _T_140 = _T_133[2:0]; // @[LZD.scala 49:59]
  assign _T_141 = _T_134 ? _T_139 : _T_140; // @[LZD.scala 49:35]
  assign _T_143 = {_T_136,_T_138,_T_141}; // @[Cat.scala 29:58]
  assign _T_144 = _T_10[15:0]; // @[LZD.scala 44:32]
  assign _T_145 = _T_144[15:8]; // @[LZD.scala 43:32]
  assign _T_146 = _T_145[7:4]; // @[LZD.scala 43:32]
  assign _T_147 = _T_146[3:2]; // @[LZD.scala 43:32]
  assign _T_148 = _T_147 != 2'h0; // @[LZD.scala 39:14]
  assign _T_149 = _T_147[1]; // @[LZD.scala 39:21]
  assign _T_150 = _T_147[0]; // @[LZD.scala 39:30]
  assign _T_151 = ~ _T_150; // @[LZD.scala 39:27]
  assign _T_152 = _T_149 | _T_151; // @[LZD.scala 39:25]
  assign _T_153 = {_T_148,_T_152}; // @[Cat.scala 29:58]
  assign _T_154 = _T_146[1:0]; // @[LZD.scala 44:32]
  assign _T_155 = _T_154 != 2'h0; // @[LZD.scala 39:14]
  assign _T_156 = _T_154[1]; // @[LZD.scala 39:21]
  assign _T_157 = _T_154[0]; // @[LZD.scala 39:30]
  assign _T_158 = ~ _T_157; // @[LZD.scala 39:27]
  assign _T_159 = _T_156 | _T_158; // @[LZD.scala 39:25]
  assign _T_160 = {_T_155,_T_159}; // @[Cat.scala 29:58]
  assign _T_161 = _T_153[1]; // @[Shift.scala 12:21]
  assign _T_162 = _T_160[1]; // @[Shift.scala 12:21]
  assign _T_163 = _T_161 | _T_162; // @[LZD.scala 49:16]
  assign _T_164 = ~ _T_162; // @[LZD.scala 49:27]
  assign _T_165 = _T_161 | _T_164; // @[LZD.scala 49:25]
  assign _T_166 = _T_153[0:0]; // @[LZD.scala 49:47]
  assign _T_167 = _T_160[0:0]; // @[LZD.scala 49:59]
  assign _T_168 = _T_161 ? _T_166 : _T_167; // @[LZD.scala 49:35]
  assign _T_170 = {_T_163,_T_165,_T_168}; // @[Cat.scala 29:58]
  assign _T_171 = _T_145[3:0]; // @[LZD.scala 44:32]
  assign _T_172 = _T_171[3:2]; // @[LZD.scala 43:32]
  assign _T_173 = _T_172 != 2'h0; // @[LZD.scala 39:14]
  assign _T_174 = _T_172[1]; // @[LZD.scala 39:21]
  assign _T_175 = _T_172[0]; // @[LZD.scala 39:30]
  assign _T_176 = ~ _T_175; // @[LZD.scala 39:27]
  assign _T_177 = _T_174 | _T_176; // @[LZD.scala 39:25]
  assign _T_178 = {_T_173,_T_177}; // @[Cat.scala 29:58]
  assign _T_179 = _T_171[1:0]; // @[LZD.scala 44:32]
  assign _T_180 = _T_179 != 2'h0; // @[LZD.scala 39:14]
  assign _T_181 = _T_179[1]; // @[LZD.scala 39:21]
  assign _T_182 = _T_179[0]; // @[LZD.scala 39:30]
  assign _T_183 = ~ _T_182; // @[LZD.scala 39:27]
  assign _T_184 = _T_181 | _T_183; // @[LZD.scala 39:25]
  assign _T_185 = {_T_180,_T_184}; // @[Cat.scala 29:58]
  assign _T_186 = _T_178[1]; // @[Shift.scala 12:21]
  assign _T_187 = _T_185[1]; // @[Shift.scala 12:21]
  assign _T_188 = _T_186 | _T_187; // @[LZD.scala 49:16]
  assign _T_189 = ~ _T_187; // @[LZD.scala 49:27]
  assign _T_190 = _T_186 | _T_189; // @[LZD.scala 49:25]
  assign _T_191 = _T_178[0:0]; // @[LZD.scala 49:47]
  assign _T_192 = _T_185[0:0]; // @[LZD.scala 49:59]
  assign _T_193 = _T_186 ? _T_191 : _T_192; // @[LZD.scala 49:35]
  assign _T_195 = {_T_188,_T_190,_T_193}; // @[Cat.scala 29:58]
  assign _T_196 = _T_170[2]; // @[Shift.scala 12:21]
  assign _T_197 = _T_195[2]; // @[Shift.scala 12:21]
  assign _T_198 = _T_196 | _T_197; // @[LZD.scala 49:16]
  assign _T_199 = ~ _T_197; // @[LZD.scala 49:27]
  assign _T_200 = _T_196 | _T_199; // @[LZD.scala 49:25]
  assign _T_201 = _T_170[1:0]; // @[LZD.scala 49:47]
  assign _T_202 = _T_195[1:0]; // @[LZD.scala 49:59]
  assign _T_203 = _T_196 ? _T_201 : _T_202; // @[LZD.scala 49:35]
  assign _T_205 = {_T_198,_T_200,_T_203}; // @[Cat.scala 29:58]
  assign _T_206 = _T_144[7:0]; // @[LZD.scala 44:32]
  assign _T_207 = _T_206[7:4]; // @[LZD.scala 43:32]
  assign _T_208 = _T_207[3:2]; // @[LZD.scala 43:32]
  assign _T_209 = _T_208 != 2'h0; // @[LZD.scala 39:14]
  assign _T_210 = _T_208[1]; // @[LZD.scala 39:21]
  assign _T_211 = _T_208[0]; // @[LZD.scala 39:30]
  assign _T_212 = ~ _T_211; // @[LZD.scala 39:27]
  assign _T_213 = _T_210 | _T_212; // @[LZD.scala 39:25]
  assign _T_214 = {_T_209,_T_213}; // @[Cat.scala 29:58]
  assign _T_215 = _T_207[1:0]; // @[LZD.scala 44:32]
  assign _T_216 = _T_215 != 2'h0; // @[LZD.scala 39:14]
  assign _T_217 = _T_215[1]; // @[LZD.scala 39:21]
  assign _T_218 = _T_215[0]; // @[LZD.scala 39:30]
  assign _T_219 = ~ _T_218; // @[LZD.scala 39:27]
  assign _T_220 = _T_217 | _T_219; // @[LZD.scala 39:25]
  assign _T_221 = {_T_216,_T_220}; // @[Cat.scala 29:58]
  assign _T_222 = _T_214[1]; // @[Shift.scala 12:21]
  assign _T_223 = _T_221[1]; // @[Shift.scala 12:21]
  assign _T_224 = _T_222 | _T_223; // @[LZD.scala 49:16]
  assign _T_225 = ~ _T_223; // @[LZD.scala 49:27]
  assign _T_226 = _T_222 | _T_225; // @[LZD.scala 49:25]
  assign _T_227 = _T_214[0:0]; // @[LZD.scala 49:47]
  assign _T_228 = _T_221[0:0]; // @[LZD.scala 49:59]
  assign _T_229 = _T_222 ? _T_227 : _T_228; // @[LZD.scala 49:35]
  assign _T_231 = {_T_224,_T_226,_T_229}; // @[Cat.scala 29:58]
  assign _T_232 = _T_206[3:0]; // @[LZD.scala 44:32]
  assign _T_233 = _T_232[3:2]; // @[LZD.scala 43:32]
  assign _T_234 = _T_233 != 2'h0; // @[LZD.scala 39:14]
  assign _T_235 = _T_233[1]; // @[LZD.scala 39:21]
  assign _T_236 = _T_233[0]; // @[LZD.scala 39:30]
  assign _T_237 = ~ _T_236; // @[LZD.scala 39:27]
  assign _T_238 = _T_235 | _T_237; // @[LZD.scala 39:25]
  assign _T_239 = {_T_234,_T_238}; // @[Cat.scala 29:58]
  assign _T_240 = _T_232[1:0]; // @[LZD.scala 44:32]
  assign _T_241 = _T_240 != 2'h0; // @[LZD.scala 39:14]
  assign _T_242 = _T_240[1]; // @[LZD.scala 39:21]
  assign _T_243 = _T_240[0]; // @[LZD.scala 39:30]
  assign _T_244 = ~ _T_243; // @[LZD.scala 39:27]
  assign _T_245 = _T_242 | _T_244; // @[LZD.scala 39:25]
  assign _T_246 = {_T_241,_T_245}; // @[Cat.scala 29:58]
  assign _T_247 = _T_239[1]; // @[Shift.scala 12:21]
  assign _T_248 = _T_246[1]; // @[Shift.scala 12:21]
  assign _T_249 = _T_247 | _T_248; // @[LZD.scala 49:16]
  assign _T_250 = ~ _T_248; // @[LZD.scala 49:27]
  assign _T_251 = _T_247 | _T_250; // @[LZD.scala 49:25]
  assign _T_252 = _T_239[0:0]; // @[LZD.scala 49:47]
  assign _T_253 = _T_246[0:0]; // @[LZD.scala 49:59]
  assign _T_254 = _T_247 ? _T_252 : _T_253; // @[LZD.scala 49:35]
  assign _T_256 = {_T_249,_T_251,_T_254}; // @[Cat.scala 29:58]
  assign _T_257 = _T_231[2]; // @[Shift.scala 12:21]
  assign _T_258 = _T_256[2]; // @[Shift.scala 12:21]
  assign _T_259 = _T_257 | _T_258; // @[LZD.scala 49:16]
  assign _T_260 = ~ _T_258; // @[LZD.scala 49:27]
  assign _T_261 = _T_257 | _T_260; // @[LZD.scala 49:25]
  assign _T_262 = _T_231[1:0]; // @[LZD.scala 49:47]
  assign _T_263 = _T_256[1:0]; // @[LZD.scala 49:59]
  assign _T_264 = _T_257 ? _T_262 : _T_263; // @[LZD.scala 49:35]
  assign _T_266 = {_T_259,_T_261,_T_264}; // @[Cat.scala 29:58]
  assign _T_267 = _T_205[3]; // @[Shift.scala 12:21]
  assign _T_268 = _T_266[3]; // @[Shift.scala 12:21]
  assign _T_269 = _T_267 | _T_268; // @[LZD.scala 49:16]
  assign _T_270 = ~ _T_268; // @[LZD.scala 49:27]
  assign _T_271 = _T_267 | _T_270; // @[LZD.scala 49:25]
  assign _T_272 = _T_205[2:0]; // @[LZD.scala 49:47]
  assign _T_273 = _T_266[2:0]; // @[LZD.scala 49:59]
  assign _T_274 = _T_267 ? _T_272 : _T_273; // @[LZD.scala 49:35]
  assign _T_276 = {_T_269,_T_271,_T_274}; // @[Cat.scala 29:58]
  assign _T_277 = _T_143[4]; // @[Shift.scala 12:21]
  assign _T_278 = _T_276[4]; // @[Shift.scala 12:21]
  assign _T_279 = _T_277 | _T_278; // @[LZD.scala 49:16]
  assign _T_280 = ~ _T_278; // @[LZD.scala 49:27]
  assign _T_281 = _T_277 | _T_280; // @[LZD.scala 49:25]
  assign _T_282 = _T_143[3:0]; // @[LZD.scala 49:47]
  assign _T_283 = _T_276[3:0]; // @[LZD.scala 49:59]
  assign _T_284 = _T_277 ? _T_282 : _T_283; // @[LZD.scala 49:35]
  assign _T_286 = {_T_279,_T_281,_T_284}; // @[Cat.scala 29:58]
  assign _T_287 = quireXOR[30:0]; // @[LZD.scala 44:32]
  assign _T_288 = _T_287[30:15]; // @[LZD.scala 43:32]
  assign _T_289 = _T_288[15:8]; // @[LZD.scala 43:32]
  assign _T_290 = _T_289[7:4]; // @[LZD.scala 43:32]
  assign _T_291 = _T_290[3:2]; // @[LZD.scala 43:32]
  assign _T_292 = _T_291 != 2'h0; // @[LZD.scala 39:14]
  assign _T_293 = _T_291[1]; // @[LZD.scala 39:21]
  assign _T_294 = _T_291[0]; // @[LZD.scala 39:30]
  assign _T_295 = ~ _T_294; // @[LZD.scala 39:27]
  assign _T_296 = _T_293 | _T_295; // @[LZD.scala 39:25]
  assign _T_297 = {_T_292,_T_296}; // @[Cat.scala 29:58]
  assign _T_298 = _T_290[1:0]; // @[LZD.scala 44:32]
  assign _T_299 = _T_298 != 2'h0; // @[LZD.scala 39:14]
  assign _T_300 = _T_298[1]; // @[LZD.scala 39:21]
  assign _T_301 = _T_298[0]; // @[LZD.scala 39:30]
  assign _T_302 = ~ _T_301; // @[LZD.scala 39:27]
  assign _T_303 = _T_300 | _T_302; // @[LZD.scala 39:25]
  assign _T_304 = {_T_299,_T_303}; // @[Cat.scala 29:58]
  assign _T_305 = _T_297[1]; // @[Shift.scala 12:21]
  assign _T_306 = _T_304[1]; // @[Shift.scala 12:21]
  assign _T_307 = _T_305 | _T_306; // @[LZD.scala 49:16]
  assign _T_308 = ~ _T_306; // @[LZD.scala 49:27]
  assign _T_309 = _T_305 | _T_308; // @[LZD.scala 49:25]
  assign _T_310 = _T_297[0:0]; // @[LZD.scala 49:47]
  assign _T_311 = _T_304[0:0]; // @[LZD.scala 49:59]
  assign _T_312 = _T_305 ? _T_310 : _T_311; // @[LZD.scala 49:35]
  assign _T_314 = {_T_307,_T_309,_T_312}; // @[Cat.scala 29:58]
  assign _T_315 = _T_289[3:0]; // @[LZD.scala 44:32]
  assign _T_316 = _T_315[3:2]; // @[LZD.scala 43:32]
  assign _T_317 = _T_316 != 2'h0; // @[LZD.scala 39:14]
  assign _T_318 = _T_316[1]; // @[LZD.scala 39:21]
  assign _T_319 = _T_316[0]; // @[LZD.scala 39:30]
  assign _T_320 = ~ _T_319; // @[LZD.scala 39:27]
  assign _T_321 = _T_318 | _T_320; // @[LZD.scala 39:25]
  assign _T_322 = {_T_317,_T_321}; // @[Cat.scala 29:58]
  assign _T_323 = _T_315[1:0]; // @[LZD.scala 44:32]
  assign _T_324 = _T_323 != 2'h0; // @[LZD.scala 39:14]
  assign _T_325 = _T_323[1]; // @[LZD.scala 39:21]
  assign _T_326 = _T_323[0]; // @[LZD.scala 39:30]
  assign _T_327 = ~ _T_326; // @[LZD.scala 39:27]
  assign _T_328 = _T_325 | _T_327; // @[LZD.scala 39:25]
  assign _T_329 = {_T_324,_T_328}; // @[Cat.scala 29:58]
  assign _T_330 = _T_322[1]; // @[Shift.scala 12:21]
  assign _T_331 = _T_329[1]; // @[Shift.scala 12:21]
  assign _T_332 = _T_330 | _T_331; // @[LZD.scala 49:16]
  assign _T_333 = ~ _T_331; // @[LZD.scala 49:27]
  assign _T_334 = _T_330 | _T_333; // @[LZD.scala 49:25]
  assign _T_335 = _T_322[0:0]; // @[LZD.scala 49:47]
  assign _T_336 = _T_329[0:0]; // @[LZD.scala 49:59]
  assign _T_337 = _T_330 ? _T_335 : _T_336; // @[LZD.scala 49:35]
  assign _T_339 = {_T_332,_T_334,_T_337}; // @[Cat.scala 29:58]
  assign _T_340 = _T_314[2]; // @[Shift.scala 12:21]
  assign _T_341 = _T_339[2]; // @[Shift.scala 12:21]
  assign _T_342 = _T_340 | _T_341; // @[LZD.scala 49:16]
  assign _T_343 = ~ _T_341; // @[LZD.scala 49:27]
  assign _T_344 = _T_340 | _T_343; // @[LZD.scala 49:25]
  assign _T_345 = _T_314[1:0]; // @[LZD.scala 49:47]
  assign _T_346 = _T_339[1:0]; // @[LZD.scala 49:59]
  assign _T_347 = _T_340 ? _T_345 : _T_346; // @[LZD.scala 49:35]
  assign _T_349 = {_T_342,_T_344,_T_347}; // @[Cat.scala 29:58]
  assign _T_350 = _T_288[7:0]; // @[LZD.scala 44:32]
  assign _T_351 = _T_350[7:4]; // @[LZD.scala 43:32]
  assign _T_352 = _T_351[3:2]; // @[LZD.scala 43:32]
  assign _T_353 = _T_352 != 2'h0; // @[LZD.scala 39:14]
  assign _T_354 = _T_352[1]; // @[LZD.scala 39:21]
  assign _T_355 = _T_352[0]; // @[LZD.scala 39:30]
  assign _T_356 = ~ _T_355; // @[LZD.scala 39:27]
  assign _T_357 = _T_354 | _T_356; // @[LZD.scala 39:25]
  assign _T_358 = {_T_353,_T_357}; // @[Cat.scala 29:58]
  assign _T_359 = _T_351[1:0]; // @[LZD.scala 44:32]
  assign _T_360 = _T_359 != 2'h0; // @[LZD.scala 39:14]
  assign _T_361 = _T_359[1]; // @[LZD.scala 39:21]
  assign _T_362 = _T_359[0]; // @[LZD.scala 39:30]
  assign _T_363 = ~ _T_362; // @[LZD.scala 39:27]
  assign _T_364 = _T_361 | _T_363; // @[LZD.scala 39:25]
  assign _T_365 = {_T_360,_T_364}; // @[Cat.scala 29:58]
  assign _T_366 = _T_358[1]; // @[Shift.scala 12:21]
  assign _T_367 = _T_365[1]; // @[Shift.scala 12:21]
  assign _T_368 = _T_366 | _T_367; // @[LZD.scala 49:16]
  assign _T_369 = ~ _T_367; // @[LZD.scala 49:27]
  assign _T_370 = _T_366 | _T_369; // @[LZD.scala 49:25]
  assign _T_371 = _T_358[0:0]; // @[LZD.scala 49:47]
  assign _T_372 = _T_365[0:0]; // @[LZD.scala 49:59]
  assign _T_373 = _T_366 ? _T_371 : _T_372; // @[LZD.scala 49:35]
  assign _T_375 = {_T_368,_T_370,_T_373}; // @[Cat.scala 29:58]
  assign _T_376 = _T_350[3:0]; // @[LZD.scala 44:32]
  assign _T_377 = _T_376[3:2]; // @[LZD.scala 43:32]
  assign _T_378 = _T_377 != 2'h0; // @[LZD.scala 39:14]
  assign _T_379 = _T_377[1]; // @[LZD.scala 39:21]
  assign _T_380 = _T_377[0]; // @[LZD.scala 39:30]
  assign _T_381 = ~ _T_380; // @[LZD.scala 39:27]
  assign _T_382 = _T_379 | _T_381; // @[LZD.scala 39:25]
  assign _T_383 = {_T_378,_T_382}; // @[Cat.scala 29:58]
  assign _T_384 = _T_376[1:0]; // @[LZD.scala 44:32]
  assign _T_385 = _T_384 != 2'h0; // @[LZD.scala 39:14]
  assign _T_386 = _T_384[1]; // @[LZD.scala 39:21]
  assign _T_387 = _T_384[0]; // @[LZD.scala 39:30]
  assign _T_388 = ~ _T_387; // @[LZD.scala 39:27]
  assign _T_389 = _T_386 | _T_388; // @[LZD.scala 39:25]
  assign _T_390 = {_T_385,_T_389}; // @[Cat.scala 29:58]
  assign _T_391 = _T_383[1]; // @[Shift.scala 12:21]
  assign _T_392 = _T_390[1]; // @[Shift.scala 12:21]
  assign _T_393 = _T_391 | _T_392; // @[LZD.scala 49:16]
  assign _T_394 = ~ _T_392; // @[LZD.scala 49:27]
  assign _T_395 = _T_391 | _T_394; // @[LZD.scala 49:25]
  assign _T_396 = _T_383[0:0]; // @[LZD.scala 49:47]
  assign _T_397 = _T_390[0:0]; // @[LZD.scala 49:59]
  assign _T_398 = _T_391 ? _T_396 : _T_397; // @[LZD.scala 49:35]
  assign _T_400 = {_T_393,_T_395,_T_398}; // @[Cat.scala 29:58]
  assign _T_401 = _T_375[2]; // @[Shift.scala 12:21]
  assign _T_402 = _T_400[2]; // @[Shift.scala 12:21]
  assign _T_403 = _T_401 | _T_402; // @[LZD.scala 49:16]
  assign _T_404 = ~ _T_402; // @[LZD.scala 49:27]
  assign _T_405 = _T_401 | _T_404; // @[LZD.scala 49:25]
  assign _T_406 = _T_375[1:0]; // @[LZD.scala 49:47]
  assign _T_407 = _T_400[1:0]; // @[LZD.scala 49:59]
  assign _T_408 = _T_401 ? _T_406 : _T_407; // @[LZD.scala 49:35]
  assign _T_410 = {_T_403,_T_405,_T_408}; // @[Cat.scala 29:58]
  assign _T_411 = _T_349[3]; // @[Shift.scala 12:21]
  assign _T_412 = _T_410[3]; // @[Shift.scala 12:21]
  assign _T_413 = _T_411 | _T_412; // @[LZD.scala 49:16]
  assign _T_414 = ~ _T_412; // @[LZD.scala 49:27]
  assign _T_415 = _T_411 | _T_414; // @[LZD.scala 49:25]
  assign _T_416 = _T_349[2:0]; // @[LZD.scala 49:47]
  assign _T_417 = _T_410[2:0]; // @[LZD.scala 49:59]
  assign _T_418 = _T_411 ? _T_416 : _T_417; // @[LZD.scala 49:35]
  assign _T_420 = {_T_413,_T_415,_T_418}; // @[Cat.scala 29:58]
  assign _T_421 = _T_287[14:0]; // @[LZD.scala 44:32]
  assign _T_422 = _T_421[14:7]; // @[LZD.scala 43:32]
  assign _T_423 = _T_422[7:4]; // @[LZD.scala 43:32]
  assign _T_424 = _T_423[3:2]; // @[LZD.scala 43:32]
  assign _T_425 = _T_424 != 2'h0; // @[LZD.scala 39:14]
  assign _T_426 = _T_424[1]; // @[LZD.scala 39:21]
  assign _T_427 = _T_424[0]; // @[LZD.scala 39:30]
  assign _T_428 = ~ _T_427; // @[LZD.scala 39:27]
  assign _T_429 = _T_426 | _T_428; // @[LZD.scala 39:25]
  assign _T_430 = {_T_425,_T_429}; // @[Cat.scala 29:58]
  assign _T_431 = _T_423[1:0]; // @[LZD.scala 44:32]
  assign _T_432 = _T_431 != 2'h0; // @[LZD.scala 39:14]
  assign _T_433 = _T_431[1]; // @[LZD.scala 39:21]
  assign _T_434 = _T_431[0]; // @[LZD.scala 39:30]
  assign _T_435 = ~ _T_434; // @[LZD.scala 39:27]
  assign _T_436 = _T_433 | _T_435; // @[LZD.scala 39:25]
  assign _T_437 = {_T_432,_T_436}; // @[Cat.scala 29:58]
  assign _T_438 = _T_430[1]; // @[Shift.scala 12:21]
  assign _T_439 = _T_437[1]; // @[Shift.scala 12:21]
  assign _T_440 = _T_438 | _T_439; // @[LZD.scala 49:16]
  assign _T_441 = ~ _T_439; // @[LZD.scala 49:27]
  assign _T_442 = _T_438 | _T_441; // @[LZD.scala 49:25]
  assign _T_443 = _T_430[0:0]; // @[LZD.scala 49:47]
  assign _T_444 = _T_437[0:0]; // @[LZD.scala 49:59]
  assign _T_445 = _T_438 ? _T_443 : _T_444; // @[LZD.scala 49:35]
  assign _T_447 = {_T_440,_T_442,_T_445}; // @[Cat.scala 29:58]
  assign _T_448 = _T_422[3:0]; // @[LZD.scala 44:32]
  assign _T_449 = _T_448[3:2]; // @[LZD.scala 43:32]
  assign _T_450 = _T_449 != 2'h0; // @[LZD.scala 39:14]
  assign _T_451 = _T_449[1]; // @[LZD.scala 39:21]
  assign _T_452 = _T_449[0]; // @[LZD.scala 39:30]
  assign _T_453 = ~ _T_452; // @[LZD.scala 39:27]
  assign _T_454 = _T_451 | _T_453; // @[LZD.scala 39:25]
  assign _T_455 = {_T_450,_T_454}; // @[Cat.scala 29:58]
  assign _T_456 = _T_448[1:0]; // @[LZD.scala 44:32]
  assign _T_457 = _T_456 != 2'h0; // @[LZD.scala 39:14]
  assign _T_458 = _T_456[1]; // @[LZD.scala 39:21]
  assign _T_459 = _T_456[0]; // @[LZD.scala 39:30]
  assign _T_460 = ~ _T_459; // @[LZD.scala 39:27]
  assign _T_461 = _T_458 | _T_460; // @[LZD.scala 39:25]
  assign _T_462 = {_T_457,_T_461}; // @[Cat.scala 29:58]
  assign _T_463 = _T_455[1]; // @[Shift.scala 12:21]
  assign _T_464 = _T_462[1]; // @[Shift.scala 12:21]
  assign _T_465 = _T_463 | _T_464; // @[LZD.scala 49:16]
  assign _T_466 = ~ _T_464; // @[LZD.scala 49:27]
  assign _T_467 = _T_463 | _T_466; // @[LZD.scala 49:25]
  assign _T_468 = _T_455[0:0]; // @[LZD.scala 49:47]
  assign _T_469 = _T_462[0:0]; // @[LZD.scala 49:59]
  assign _T_470 = _T_463 ? _T_468 : _T_469; // @[LZD.scala 49:35]
  assign _T_472 = {_T_465,_T_467,_T_470}; // @[Cat.scala 29:58]
  assign _T_473 = _T_447[2]; // @[Shift.scala 12:21]
  assign _T_474 = _T_472[2]; // @[Shift.scala 12:21]
  assign _T_475 = _T_473 | _T_474; // @[LZD.scala 49:16]
  assign _T_476 = ~ _T_474; // @[LZD.scala 49:27]
  assign _T_477 = _T_473 | _T_476; // @[LZD.scala 49:25]
  assign _T_478 = _T_447[1:0]; // @[LZD.scala 49:47]
  assign _T_479 = _T_472[1:0]; // @[LZD.scala 49:59]
  assign _T_480 = _T_473 ? _T_478 : _T_479; // @[LZD.scala 49:35]
  assign _T_482 = {_T_475,_T_477,_T_480}; // @[Cat.scala 29:58]
  assign _T_483 = _T_421[6:0]; // @[LZD.scala 44:32]
  assign _T_484 = _T_483[6:3]; // @[LZD.scala 43:32]
  assign _T_485 = _T_484[3:2]; // @[LZD.scala 43:32]
  assign _T_486 = _T_485 != 2'h0; // @[LZD.scala 39:14]
  assign _T_487 = _T_485[1]; // @[LZD.scala 39:21]
  assign _T_488 = _T_485[0]; // @[LZD.scala 39:30]
  assign _T_489 = ~ _T_488; // @[LZD.scala 39:27]
  assign _T_490 = _T_487 | _T_489; // @[LZD.scala 39:25]
  assign _T_491 = {_T_486,_T_490}; // @[Cat.scala 29:58]
  assign _T_492 = _T_484[1:0]; // @[LZD.scala 44:32]
  assign _T_493 = _T_492 != 2'h0; // @[LZD.scala 39:14]
  assign _T_494 = _T_492[1]; // @[LZD.scala 39:21]
  assign _T_495 = _T_492[0]; // @[LZD.scala 39:30]
  assign _T_496 = ~ _T_495; // @[LZD.scala 39:27]
  assign _T_497 = _T_494 | _T_496; // @[LZD.scala 39:25]
  assign _T_498 = {_T_493,_T_497}; // @[Cat.scala 29:58]
  assign _T_499 = _T_491[1]; // @[Shift.scala 12:21]
  assign _T_500 = _T_498[1]; // @[Shift.scala 12:21]
  assign _T_501 = _T_499 | _T_500; // @[LZD.scala 49:16]
  assign _T_502 = ~ _T_500; // @[LZD.scala 49:27]
  assign _T_503 = _T_499 | _T_502; // @[LZD.scala 49:25]
  assign _T_504 = _T_491[0:0]; // @[LZD.scala 49:47]
  assign _T_505 = _T_498[0:0]; // @[LZD.scala 49:59]
  assign _T_506 = _T_499 ? _T_504 : _T_505; // @[LZD.scala 49:35]
  assign _T_508 = {_T_501,_T_503,_T_506}; // @[Cat.scala 29:58]
  assign _T_509 = _T_483[2:0]; // @[LZD.scala 44:32]
  assign _T_510 = _T_509[2:1]; // @[LZD.scala 43:32]
  assign _T_511 = _T_510 != 2'h0; // @[LZD.scala 39:14]
  assign _T_512 = _T_510[1]; // @[LZD.scala 39:21]
  assign _T_513 = _T_510[0]; // @[LZD.scala 39:30]
  assign _T_514 = ~ _T_513; // @[LZD.scala 39:27]
  assign _T_515 = _T_512 | _T_514; // @[LZD.scala 39:25]
  assign _T_516 = {_T_511,_T_515}; // @[Cat.scala 29:58]
  assign _T_517 = _T_509[0:0]; // @[LZD.scala 44:32]
  assign _T_519 = _T_516[1]; // @[Shift.scala 12:21]
  assign _T_521 = _T_516[0:0]; // @[LZD.scala 55:32]
  assign _T_522 = _T_519 ? _T_521 : _T_517; // @[LZD.scala 55:20]
  assign _T_523 = {_T_519,_T_522}; // @[Cat.scala 29:58]
  assign _T_524 = _T_508[2]; // @[Shift.scala 12:21]
  assign _T_526 = _T_508[1:0]; // @[LZD.scala 55:32]
  assign _T_527 = _T_524 ? _T_526 : _T_523; // @[LZD.scala 55:20]
  assign _T_528 = {_T_524,_T_527}; // @[Cat.scala 29:58]
  assign _T_529 = _T_482[3]; // @[Shift.scala 12:21]
  assign _T_531 = _T_482[2:0]; // @[LZD.scala 55:32]
  assign _T_532 = _T_529 ? _T_531 : _T_528; // @[LZD.scala 55:20]
  assign _T_533 = {_T_529,_T_532}; // @[Cat.scala 29:58]
  assign _T_534 = _T_420[4]; // @[Shift.scala 12:21]
  assign _T_536 = _T_420[3:0]; // @[LZD.scala 55:32]
  assign _T_537 = _T_534 ? _T_536 : _T_533; // @[LZD.scala 55:20]
  assign _T_538 = {_T_534,_T_537}; // @[Cat.scala 29:58]
  assign _T_539 = _T_286[5]; // @[Shift.scala 12:21]
  assign _T_541 = _T_286[4:0]; // @[LZD.scala 55:32]
  assign _T_542 = _T_539 ? _T_541 : _T_538; // @[LZD.scala 55:20]
  assign scaleBias = {1'h1,_T_539,_T_542}; // @[Cat.scala 29:58]
  assign _T_543 = $signed(scaleBias); // @[QuireToPosit.scala 61:53]
  assign _GEN_2 = {{1{_T_543[6]}},_T_543}; // @[QuireToPosit.scala 61:41]
  assign _T_545 = $signed(8'sh27) + $signed(_GEN_2); // @[QuireToPosit.scala 61:41]
  assign realScale = $signed(_T_545); // @[QuireToPosit.scala 61:41]
  assign underflow = $signed(realScale) < $signed(-8'shd); // @[QuireToPosit.scala 62:41]
  assign overflow = $signed(realScale) > $signed(8'shc); // @[QuireToPosit.scala 63:35]
  assign _T_546 = underflow ? $signed(-8'shd) : $signed(realScale); // @[Mux.scala 87:16]
  assign _T_547 = overflow ? $signed(8'shc) : $signed(_T_546); // @[Mux.scala 87:16]
  assign _T_548 = realScale[7:7]; // @[Abs.scala 10:21]
  assign _T_550 = _T_548 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_551 = $unsigned(realScale); // @[Abs.scala 10:31]
  assign _T_552 = _T_550 ^ _T_551; // @[Abs.scala 10:26]
  assign _GEN_3 = {{7'd0}, _T_548}; // @[Abs.scala 10:39]
  assign absRealScale = _T_552 + _GEN_3; // @[Abs.scala 10:39]
  assign _T_555 = absRealScale < 8'h40; // @[Shift.scala 16:24]
  assign _T_556 = absRealScale[5:0]; // @[Shift.scala 17:37]
  assign _T_557 = _T_556[5]; // @[Shift.scala 12:21]
  assign _T_558 = io_quireIn[31:0]; // @[Shift.scala 64:52]
  assign _T_560 = {_T_558,32'h0}; // @[Cat.scala 29:58]
  assign _T_561 = _T_557 ? _T_560 : io_quireIn; // @[Shift.scala 64:27]
  assign _T_562 = _T_556[4:0]; // @[Shift.scala 66:70]
  assign _T_563 = _T_562[4]; // @[Shift.scala 12:21]
  assign _T_564 = _T_561[47:0]; // @[Shift.scala 64:52]
  assign _T_566 = {_T_564,16'h0}; // @[Cat.scala 29:58]
  assign _T_567 = _T_563 ? _T_566 : _T_561; // @[Shift.scala 64:27]
  assign _T_568 = _T_562[3:0]; // @[Shift.scala 66:70]
  assign _T_569 = _T_568[3]; // @[Shift.scala 12:21]
  assign _T_570 = _T_567[55:0]; // @[Shift.scala 64:52]
  assign _T_572 = {_T_570,8'h0}; // @[Cat.scala 29:58]
  assign _T_573 = _T_569 ? _T_572 : _T_567; // @[Shift.scala 64:27]
  assign _T_574 = _T_568[2:0]; // @[Shift.scala 66:70]
  assign _T_575 = _T_574[2]; // @[Shift.scala 12:21]
  assign _T_576 = _T_573[59:0]; // @[Shift.scala 64:52]
  assign _T_578 = {_T_576,4'h0}; // @[Cat.scala 29:58]
  assign _T_579 = _T_575 ? _T_578 : _T_573; // @[Shift.scala 64:27]
  assign _T_580 = _T_574[1:0]; // @[Shift.scala 66:70]
  assign _T_581 = _T_580[1]; // @[Shift.scala 12:21]
  assign _T_582 = _T_579[61:0]; // @[Shift.scala 64:52]
  assign _T_584 = {_T_582,2'h0}; // @[Cat.scala 29:58]
  assign _T_585 = _T_581 ? _T_584 : _T_579; // @[Shift.scala 64:27]
  assign _T_586 = _T_580[0:0]; // @[Shift.scala 66:70]
  assign _T_588 = _T_585[62:0]; // @[Shift.scala 64:52]
  assign _T_589 = {_T_588,1'h0}; // @[Cat.scala 29:58]
  assign _T_590 = _T_586 ? _T_589 : _T_585; // @[Shift.scala 64:27]
  assign quireLeftShift = _T_555 ? _T_590 : 64'h0; // @[Shift.scala 16:10]
  assign _T_595 = io_quireIn[63:32]; // @[Shift.scala 77:66]
  assign _T_596 = {32'h0,_T_595}; // @[Cat.scala 29:58]
  assign _T_597 = _T_557 ? _T_596 : io_quireIn; // @[Shift.scala 77:22]
  assign _T_601 = _T_597[63:16]; // @[Shift.scala 77:66]
  assign _T_602 = {16'h0,_T_601}; // @[Cat.scala 29:58]
  assign _T_603 = _T_563 ? _T_602 : _T_597; // @[Shift.scala 77:22]
  assign _T_607 = _T_603[63:8]; // @[Shift.scala 77:66]
  assign _T_608 = {8'h0,_T_607}; // @[Cat.scala 29:58]
  assign _T_609 = _T_569 ? _T_608 : _T_603; // @[Shift.scala 77:22]
  assign _T_613 = _T_609[63:4]; // @[Shift.scala 77:66]
  assign _T_614 = {4'h0,_T_613}; // @[Cat.scala 29:58]
  assign _T_615 = _T_575 ? _T_614 : _T_609; // @[Shift.scala 77:22]
  assign _T_619 = _T_615[63:2]; // @[Shift.scala 77:66]
  assign _T_620 = {2'h0,_T_619}; // @[Cat.scala 29:58]
  assign _T_621 = _T_581 ? _T_620 : _T_615; // @[Shift.scala 77:22]
  assign _T_624 = _T_621[63:1]; // @[Shift.scala 77:66]
  assign _T_625 = {1'h0,_T_624}; // @[Cat.scala 29:58]
  assign _T_626 = _T_586 ? _T_625 : _T_621; // @[Shift.scala 77:22]
  assign quireRightShift = _T_555 ? _T_626 : 64'h0; // @[Shift.scala 27:10]
  assign _T_628 = quireLeftShift[23:18]; // @[QuireToPosit.scala 89:49]
  assign _T_629 = quireLeftShift[17:0]; // @[QuireToPosit.scala 90:127]
  assign _T_630 = _T_629 != 18'h0; // @[QuireToPosit.scala 90:154]
  assign realFGRSTmp1 = {_T_628,_T_630}; // @[Cat.scala 29:58]
  assign _T_631 = quireRightShift[23:18]; // @[QuireToPosit.scala 91:50]
  assign _T_632 = quireRightShift[17:0]; // @[QuireToPosit.scala 92:128]
  assign _T_633 = _T_632 != 18'h0; // @[QuireToPosit.scala 92:155]
  assign realFGRSTmp2 = {_T_631,_T_633}; // @[Cat.scala 29:58]
  assign realFGRS = _T_548 ? realFGRSTmp1 : realFGRSTmp2; // @[QuireToPosit.scala 93:34]
  assign outRawFloat_fraction = realFGRS[6:3]; // @[QuireToPosit.scala 95:46]
  assign outRawFloat_grs = realFGRS[2:0]; // @[QuireToPosit.scala 96:46]
  assign _GEN_4 = _T_547[4:0]; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  assign outRawFloat_scale = $signed(_GEN_4); // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  assign _T_638 = outRawFloat_scale[0]; // @[convert.scala 46:61]
  assign _T_639 = ~ _T_638; // @[convert.scala 46:52]
  assign _T_641 = _T_2 ? _T_639 : _T_638; // @[convert.scala 46:42]
  assign _T_642 = outRawFloat_scale[4:1]; // @[convert.scala 48:34]
  assign _T_643 = _T_642[3:3]; // @[convert.scala 49:36]
  assign _T_645 = ~ _T_642; // @[convert.scala 50:36]
  assign _T_646 = $signed(_T_645); // @[convert.scala 50:36]
  assign _T_647 = _T_643 ? $signed(_T_646) : $signed(_T_642); // @[convert.scala 50:28]
  assign _T_648 = _T_643 ^ _T_2; // @[convert.scala 51:31]
  assign _T_649 = ~ _T_648; // @[convert.scala 52:43]
  assign _T_653 = {_T_649,_T_648,_T_641,outRawFloat_fraction,outRawFloat_grs}; // @[Cat.scala 29:58]
  assign _T_654 = $unsigned(_T_647); // @[Shift.scala 39:17]
  assign _T_655 = _T_654 < 4'ha; // @[Shift.scala 39:24]
  assign _T_657 = _T_653[9:8]; // @[Shift.scala 90:30]
  assign _T_658 = _T_653[7:0]; // @[Shift.scala 90:48]
  assign _T_659 = _T_658 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{1'd0}, _T_659}; // @[Shift.scala 90:39]
  assign _T_660 = _T_657 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_661 = _T_654[3]; // @[Shift.scala 12:21]
  assign _T_662 = _T_653[9]; // @[Shift.scala 12:21]
  assign _T_664 = _T_662 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_665 = {_T_664,_T_660}; // @[Cat.scala 29:58]
  assign _T_666 = _T_661 ? _T_665 : _T_653; // @[Shift.scala 91:22]
  assign _T_667 = _T_654[2:0]; // @[Shift.scala 92:77]
  assign _T_668 = _T_666[9:4]; // @[Shift.scala 90:30]
  assign _T_669 = _T_666[3:0]; // @[Shift.scala 90:48]
  assign _T_670 = _T_669 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{5'd0}, _T_670}; // @[Shift.scala 90:39]
  assign _T_671 = _T_668 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_672 = _T_667[2]; // @[Shift.scala 12:21]
  assign _T_673 = _T_666[9]; // @[Shift.scala 12:21]
  assign _T_675 = _T_673 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_676 = {_T_675,_T_671}; // @[Cat.scala 29:58]
  assign _T_677 = _T_672 ? _T_676 : _T_666; // @[Shift.scala 91:22]
  assign _T_678 = _T_667[1:0]; // @[Shift.scala 92:77]
  assign _T_679 = _T_677[9:2]; // @[Shift.scala 90:30]
  assign _T_680 = _T_677[1:0]; // @[Shift.scala 90:48]
  assign _T_681 = _T_680 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{7'd0}, _T_681}; // @[Shift.scala 90:39]
  assign _T_682 = _T_679 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_683 = _T_678[1]; // @[Shift.scala 12:21]
  assign _T_684 = _T_677[9]; // @[Shift.scala 12:21]
  assign _T_686 = _T_684 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_687 = {_T_686,_T_682}; // @[Cat.scala 29:58]
  assign _T_688 = _T_683 ? _T_687 : _T_677; // @[Shift.scala 91:22]
  assign _T_689 = _T_678[0:0]; // @[Shift.scala 92:77]
  assign _T_690 = _T_688[9:1]; // @[Shift.scala 90:30]
  assign _T_691 = _T_688[0:0]; // @[Shift.scala 90:48]
  assign _GEN_8 = {{8'd0}, _T_691}; // @[Shift.scala 90:39]
  assign _T_693 = _T_690 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_695 = _T_688[9]; // @[Shift.scala 12:21]
  assign _T_696 = {_T_695,_T_693}; // @[Cat.scala 29:58]
  assign _T_697 = _T_689 ? _T_696 : _T_688; // @[Shift.scala 91:22]
  assign _T_700 = _T_662 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_701 = _T_655 ? _T_697 : _T_700; // @[Shift.scala 39:10]
  assign _T_702 = _T_701[3]; // @[convert.scala 55:31]
  assign _T_703 = _T_701[2]; // @[convert.scala 56:31]
  assign _T_704 = _T_701[1]; // @[convert.scala 57:31]
  assign _T_705 = _T_701[0]; // @[convert.scala 58:31]
  assign _T_706 = _T_701[9:3]; // @[convert.scala 59:69]
  assign _T_707 = _T_706 != 7'h0; // @[convert.scala 59:81]
  assign _T_708 = ~ _T_707; // @[convert.scala 59:50]
  assign _T_710 = _T_706 == 7'h7f; // @[convert.scala 60:81]
  assign _T_711 = _T_702 | _T_704; // @[convert.scala 61:44]
  assign _T_712 = _T_711 | _T_705; // @[convert.scala 61:52]
  assign _T_713 = _T_703 & _T_712; // @[convert.scala 61:36]
  assign _T_714 = ~ _T_710; // @[convert.scala 62:63]
  assign _T_715 = _T_714 & _T_713; // @[convert.scala 62:103]
  assign _T_716 = _T_708 | _T_715; // @[convert.scala 62:60]
  assign _GEN_9 = {{6'd0}, _T_716}; // @[convert.scala 63:56]
  assign _T_719 = _T_706 + _GEN_9; // @[convert.scala 63:56]
  assign _T_720 = {_T_2,_T_719}; // @[Cat.scala 29:58]
  assign io_positOut = _T_728; // @[QuireToPosit.scala 101:15]
  assign io_outValid = _T_724; // @[QuireToPosit.scala 100:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_724 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_728 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_724 <= 1'h0;
    end else begin
      _T_724 <= io_inValid;
    end
    if (io_inValid) begin
      if (outRawFloat_isNaR) begin
        _T_728 <= 8'h80;
      end else begin
        if (outRawFloat_isZero) begin
          _T_728 <= 8'h0;
        end else begin
          _T_728 <= _T_720;
        end
      end
    end
  end
endmodule
