module FMAEnc8_1(
  input         clock,
  input         reset,
  input         io_inValid_phase2,
  input  [11:0] io_signSumSig,
  input         io_sumSign,
  input  [4:0]  io_greaterScale,
  input         io_outIsNaR_phase2,
  output [7:0]  io_F,
  output        io_outValid
);
  wire [10:0] _T; // @[FMAEnc.scala 35:36]
  wire [10:0] _T_1; // @[FMAEnc.scala 35:74]
  wire [10:0] sumXor; // @[FMAEnc.scala 35:54]
  wire [7:0] _T_2; // @[LZD.scala 43:32]
  wire [3:0] _T_3; // @[LZD.scala 43:32]
  wire [1:0] _T_4; // @[LZD.scala 43:32]
  wire  _T_5; // @[LZD.scala 39:14]
  wire  _T_6; // @[LZD.scala 39:21]
  wire  _T_7; // @[LZD.scala 39:30]
  wire  _T_8; // @[LZD.scala 39:27]
  wire  _T_9; // @[LZD.scala 39:25]
  wire [1:0] _T_10; // @[Cat.scala 29:58]
  wire [1:0] _T_11; // @[LZD.scala 44:32]
  wire  _T_12; // @[LZD.scala 39:14]
  wire  _T_13; // @[LZD.scala 39:21]
  wire  _T_14; // @[LZD.scala 39:30]
  wire  _T_15; // @[LZD.scala 39:27]
  wire  _T_16; // @[LZD.scala 39:25]
  wire [1:0] _T_17; // @[Cat.scala 29:58]
  wire  _T_18; // @[Shift.scala 12:21]
  wire  _T_19; // @[Shift.scala 12:21]
  wire  _T_20; // @[LZD.scala 49:16]
  wire  _T_21; // @[LZD.scala 49:27]
  wire  _T_22; // @[LZD.scala 49:25]
  wire  _T_23; // @[LZD.scala 49:47]
  wire  _T_24; // @[LZD.scala 49:59]
  wire  _T_25; // @[LZD.scala 49:35]
  wire [2:0] _T_27; // @[Cat.scala 29:58]
  wire [3:0] _T_28; // @[LZD.scala 44:32]
  wire [1:0] _T_29; // @[LZD.scala 43:32]
  wire  _T_30; // @[LZD.scala 39:14]
  wire  _T_31; // @[LZD.scala 39:21]
  wire  _T_32; // @[LZD.scala 39:30]
  wire  _T_33; // @[LZD.scala 39:27]
  wire  _T_34; // @[LZD.scala 39:25]
  wire [1:0] _T_35; // @[Cat.scala 29:58]
  wire [1:0] _T_36; // @[LZD.scala 44:32]
  wire  _T_37; // @[LZD.scala 39:14]
  wire  _T_38; // @[LZD.scala 39:21]
  wire  _T_39; // @[LZD.scala 39:30]
  wire  _T_40; // @[LZD.scala 39:27]
  wire  _T_41; // @[LZD.scala 39:25]
  wire [1:0] _T_42; // @[Cat.scala 29:58]
  wire  _T_43; // @[Shift.scala 12:21]
  wire  _T_44; // @[Shift.scala 12:21]
  wire  _T_45; // @[LZD.scala 49:16]
  wire  _T_46; // @[LZD.scala 49:27]
  wire  _T_47; // @[LZD.scala 49:25]
  wire  _T_48; // @[LZD.scala 49:47]
  wire  _T_49; // @[LZD.scala 49:59]
  wire  _T_50; // @[LZD.scala 49:35]
  wire [2:0] _T_52; // @[Cat.scala 29:58]
  wire  _T_53; // @[Shift.scala 12:21]
  wire  _T_54; // @[Shift.scala 12:21]
  wire  _T_55; // @[LZD.scala 49:16]
  wire  _T_56; // @[LZD.scala 49:27]
  wire  _T_57; // @[LZD.scala 49:25]
  wire [1:0] _T_58; // @[LZD.scala 49:47]
  wire [1:0] _T_59; // @[LZD.scala 49:59]
  wire [1:0] _T_60; // @[LZD.scala 49:35]
  wire [3:0] _T_62; // @[Cat.scala 29:58]
  wire [2:0] _T_63; // @[LZD.scala 44:32]
  wire [1:0] _T_64; // @[LZD.scala 43:32]
  wire  _T_65; // @[LZD.scala 39:14]
  wire  _T_66; // @[LZD.scala 39:21]
  wire  _T_67; // @[LZD.scala 39:30]
  wire  _T_68; // @[LZD.scala 39:27]
  wire  _T_69; // @[LZD.scala 39:25]
  wire [1:0] _T_70; // @[Cat.scala 29:58]
  wire  _T_71; // @[LZD.scala 44:32]
  wire  _T_73; // @[Shift.scala 12:21]
  wire  _T_75; // @[LZD.scala 55:32]
  wire  _T_76; // @[LZD.scala 55:20]
  wire  _T_78; // @[Shift.scala 12:21]
  wire [2:0] _T_80; // @[Cat.scala 29:58]
  wire [2:0] _T_81; // @[LZD.scala 55:32]
  wire [2:0] _T_82; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [3:0] shiftValue; // @[FMAEnc.scala 37:24]
  wire [9:0] _T_83; // @[FMAEnc.scala 38:41]
  wire  _T_84; // @[Shift.scala 16:24]
  wire  _T_86; // @[Shift.scala 12:21]
  wire [1:0] _T_87; // @[Shift.scala 64:52]
  wire [9:0] _T_89; // @[Cat.scala 29:58]
  wire [9:0] _T_90; // @[Shift.scala 64:27]
  wire [2:0] _T_91; // @[Shift.scala 66:70]
  wire  _T_92; // @[Shift.scala 12:21]
  wire [5:0] _T_93; // @[Shift.scala 64:52]
  wire [9:0] _T_95; // @[Cat.scala 29:58]
  wire [9:0] _T_96; // @[Shift.scala 64:27]
  wire [1:0] _T_97; // @[Shift.scala 66:70]
  wire  _T_98; // @[Shift.scala 12:21]
  wire [7:0] _T_99; // @[Shift.scala 64:52]
  wire [9:0] _T_101; // @[Cat.scala 29:58]
  wire [9:0] _T_102; // @[Shift.scala 64:27]
  wire  _T_103; // @[Shift.scala 66:70]
  wire [8:0] _T_105; // @[Shift.scala 64:52]
  wire [9:0] _T_106; // @[Cat.scala 29:58]
  wire [9:0] _T_107; // @[Shift.scala 64:27]
  wire [9:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [4:0] _T_109; // @[FMAEnc.scala 41:39]
  wire [4:0] _T_110; // @[FMAEnc.scala 41:39]
  wire [4:0] _T_111; // @[Cat.scala 29:58]
  wire [4:0] _T_112; // @[FMAEnc.scala 41:64]
  wire [4:0] _T_114; // @[FMAEnc.scala 41:45]
  wire [4:0] sumScale; // @[FMAEnc.scala 41:45]
  wire [3:0] sumFrac; // @[FMAEnc.scala 42:41]
  wire [5:0] grsTmp; // @[FMAEnc.scala 45:41]
  wire [1:0] _T_115; // @[FMAEnc.scala 48:40]
  wire [3:0] _T_116; // @[FMAEnc.scala 48:56]
  wire  _T_117; // @[FMAEnc.scala 48:60]
  wire  underflow; // @[FMAEnc.scala 55:32]
  wire  overflow; // @[FMAEnc.scala 56:32]
  wire  _T_118; // @[FMAEnc.scala 65:35]
  wire  decF_isZero; // @[FMAEnc.scala 65:20]
  wire [4:0] _T_120; // @[Mux.scala 87:16]
  wire [4:0] decF_scale; // @[Mux.scala 87:16]
  wire  _T_122; // @[convert.scala 46:61]
  wire  _T_123; // @[convert.scala 46:52]
  wire  _T_125; // @[convert.scala 46:42]
  wire [3:0] _T_126; // @[convert.scala 48:34]
  wire  _T_127; // @[convert.scala 49:36]
  wire [3:0] _T_129; // @[convert.scala 50:36]
  wire [3:0] _T_130; // @[convert.scala 50:36]
  wire [3:0] _T_131; // @[convert.scala 50:28]
  wire  _T_132; // @[convert.scala 51:31]
  wire  _T_133; // @[convert.scala 52:43]
  wire [9:0] _T_137; // @[Cat.scala 29:58]
  wire [3:0] _T_138; // @[Shift.scala 39:17]
  wire  _T_139; // @[Shift.scala 39:24]
  wire [1:0] _T_141; // @[Shift.scala 90:30]
  wire [7:0] _T_142; // @[Shift.scala 90:48]
  wire  _T_143; // @[Shift.scala 90:57]
  wire [1:0] _GEN_2; // @[Shift.scala 90:39]
  wire [1:0] _T_144; // @[Shift.scala 90:39]
  wire  _T_145; // @[Shift.scala 12:21]
  wire  _T_146; // @[Shift.scala 12:21]
  wire [7:0] _T_148; // @[Bitwise.scala 71:12]
  wire [9:0] _T_149; // @[Cat.scala 29:58]
  wire [9:0] _T_150; // @[Shift.scala 91:22]
  wire [2:0] _T_151; // @[Shift.scala 92:77]
  wire [5:0] _T_152; // @[Shift.scala 90:30]
  wire [3:0] _T_153; // @[Shift.scala 90:48]
  wire  _T_154; // @[Shift.scala 90:57]
  wire [5:0] _GEN_3; // @[Shift.scala 90:39]
  wire [5:0] _T_155; // @[Shift.scala 90:39]
  wire  _T_156; // @[Shift.scala 12:21]
  wire  _T_157; // @[Shift.scala 12:21]
  wire [3:0] _T_159; // @[Bitwise.scala 71:12]
  wire [9:0] _T_160; // @[Cat.scala 29:58]
  wire [9:0] _T_161; // @[Shift.scala 91:22]
  wire [1:0] _T_162; // @[Shift.scala 92:77]
  wire [7:0] _T_163; // @[Shift.scala 90:30]
  wire [1:0] _T_164; // @[Shift.scala 90:48]
  wire  _T_165; // @[Shift.scala 90:57]
  wire [7:0] _GEN_4; // @[Shift.scala 90:39]
  wire [7:0] _T_166; // @[Shift.scala 90:39]
  wire  _T_167; // @[Shift.scala 12:21]
  wire  _T_168; // @[Shift.scala 12:21]
  wire [1:0] _T_170; // @[Bitwise.scala 71:12]
  wire [9:0] _T_171; // @[Cat.scala 29:58]
  wire [9:0] _T_172; // @[Shift.scala 91:22]
  wire  _T_173; // @[Shift.scala 92:77]
  wire [8:0] _T_174; // @[Shift.scala 90:30]
  wire  _T_175; // @[Shift.scala 90:48]
  wire [8:0] _GEN_5; // @[Shift.scala 90:39]
  wire [8:0] _T_177; // @[Shift.scala 90:39]
  wire  _T_179; // @[Shift.scala 12:21]
  wire [9:0] _T_180; // @[Cat.scala 29:58]
  wire [9:0] _T_181; // @[Shift.scala 91:22]
  wire [9:0] _T_184; // @[Bitwise.scala 71:12]
  wire [9:0] _T_185; // @[Shift.scala 39:10]
  wire  _T_186; // @[convert.scala 55:31]
  wire  _T_187; // @[convert.scala 56:31]
  wire  _T_188; // @[convert.scala 57:31]
  wire  _T_189; // @[convert.scala 58:31]
  wire [6:0] _T_190; // @[convert.scala 59:69]
  wire  _T_191; // @[convert.scala 59:81]
  wire  _T_192; // @[convert.scala 59:50]
  wire  _T_194; // @[convert.scala 60:81]
  wire  _T_195; // @[convert.scala 61:44]
  wire  _T_196; // @[convert.scala 61:52]
  wire  _T_197; // @[convert.scala 61:36]
  wire  _T_198; // @[convert.scala 62:63]
  wire  _T_199; // @[convert.scala 62:103]
  wire  _T_200; // @[convert.scala 62:60]
  wire [6:0] _GEN_6; // @[convert.scala 63:56]
  wire [6:0] _T_203; // @[convert.scala 63:56]
  wire [7:0] _T_204; // @[Cat.scala 29:58]
  reg  _T_208; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [7:0] _T_212; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  assign _T = io_signSumSig[11:1]; // @[FMAEnc.scala 35:36]
  assign _T_1 = io_signSumSig[10:0]; // @[FMAEnc.scala 35:74]
  assign sumXor = _T ^ _T_1; // @[FMAEnc.scala 35:54]
  assign _T_2 = sumXor[10:3]; // @[LZD.scala 43:32]
  assign _T_3 = _T_2[7:4]; // @[LZD.scala 43:32]
  assign _T_4 = _T_3[3:2]; // @[LZD.scala 43:32]
  assign _T_5 = _T_4 != 2'h0; // @[LZD.scala 39:14]
  assign _T_6 = _T_4[1]; // @[LZD.scala 39:21]
  assign _T_7 = _T_4[0]; // @[LZD.scala 39:30]
  assign _T_8 = ~ _T_7; // @[LZD.scala 39:27]
  assign _T_9 = _T_6 | _T_8; // @[LZD.scala 39:25]
  assign _T_10 = {_T_5,_T_9}; // @[Cat.scala 29:58]
  assign _T_11 = _T_3[1:0]; // @[LZD.scala 44:32]
  assign _T_12 = _T_11 != 2'h0; // @[LZD.scala 39:14]
  assign _T_13 = _T_11[1]; // @[LZD.scala 39:21]
  assign _T_14 = _T_11[0]; // @[LZD.scala 39:30]
  assign _T_15 = ~ _T_14; // @[LZD.scala 39:27]
  assign _T_16 = _T_13 | _T_15; // @[LZD.scala 39:25]
  assign _T_17 = {_T_12,_T_16}; // @[Cat.scala 29:58]
  assign _T_18 = _T_10[1]; // @[Shift.scala 12:21]
  assign _T_19 = _T_17[1]; // @[Shift.scala 12:21]
  assign _T_20 = _T_18 | _T_19; // @[LZD.scala 49:16]
  assign _T_21 = ~ _T_19; // @[LZD.scala 49:27]
  assign _T_22 = _T_18 | _T_21; // @[LZD.scala 49:25]
  assign _T_23 = _T_10[0:0]; // @[LZD.scala 49:47]
  assign _T_24 = _T_17[0:0]; // @[LZD.scala 49:59]
  assign _T_25 = _T_18 ? _T_23 : _T_24; // @[LZD.scala 49:35]
  assign _T_27 = {_T_20,_T_22,_T_25}; // @[Cat.scala 29:58]
  assign _T_28 = _T_2[3:0]; // @[LZD.scala 44:32]
  assign _T_29 = _T_28[3:2]; // @[LZD.scala 43:32]
  assign _T_30 = _T_29 != 2'h0; // @[LZD.scala 39:14]
  assign _T_31 = _T_29[1]; // @[LZD.scala 39:21]
  assign _T_32 = _T_29[0]; // @[LZD.scala 39:30]
  assign _T_33 = ~ _T_32; // @[LZD.scala 39:27]
  assign _T_34 = _T_31 | _T_33; // @[LZD.scala 39:25]
  assign _T_35 = {_T_30,_T_34}; // @[Cat.scala 29:58]
  assign _T_36 = _T_28[1:0]; // @[LZD.scala 44:32]
  assign _T_37 = _T_36 != 2'h0; // @[LZD.scala 39:14]
  assign _T_38 = _T_36[1]; // @[LZD.scala 39:21]
  assign _T_39 = _T_36[0]; // @[LZD.scala 39:30]
  assign _T_40 = ~ _T_39; // @[LZD.scala 39:27]
  assign _T_41 = _T_38 | _T_40; // @[LZD.scala 39:25]
  assign _T_42 = {_T_37,_T_41}; // @[Cat.scala 29:58]
  assign _T_43 = _T_35[1]; // @[Shift.scala 12:21]
  assign _T_44 = _T_42[1]; // @[Shift.scala 12:21]
  assign _T_45 = _T_43 | _T_44; // @[LZD.scala 49:16]
  assign _T_46 = ~ _T_44; // @[LZD.scala 49:27]
  assign _T_47 = _T_43 | _T_46; // @[LZD.scala 49:25]
  assign _T_48 = _T_35[0:0]; // @[LZD.scala 49:47]
  assign _T_49 = _T_42[0:0]; // @[LZD.scala 49:59]
  assign _T_50 = _T_43 ? _T_48 : _T_49; // @[LZD.scala 49:35]
  assign _T_52 = {_T_45,_T_47,_T_50}; // @[Cat.scala 29:58]
  assign _T_53 = _T_27[2]; // @[Shift.scala 12:21]
  assign _T_54 = _T_52[2]; // @[Shift.scala 12:21]
  assign _T_55 = _T_53 | _T_54; // @[LZD.scala 49:16]
  assign _T_56 = ~ _T_54; // @[LZD.scala 49:27]
  assign _T_57 = _T_53 | _T_56; // @[LZD.scala 49:25]
  assign _T_58 = _T_27[1:0]; // @[LZD.scala 49:47]
  assign _T_59 = _T_52[1:0]; // @[LZD.scala 49:59]
  assign _T_60 = _T_53 ? _T_58 : _T_59; // @[LZD.scala 49:35]
  assign _T_62 = {_T_55,_T_57,_T_60}; // @[Cat.scala 29:58]
  assign _T_63 = sumXor[2:0]; // @[LZD.scala 44:32]
  assign _T_64 = _T_63[2:1]; // @[LZD.scala 43:32]
  assign _T_65 = _T_64 != 2'h0; // @[LZD.scala 39:14]
  assign _T_66 = _T_64[1]; // @[LZD.scala 39:21]
  assign _T_67 = _T_64[0]; // @[LZD.scala 39:30]
  assign _T_68 = ~ _T_67; // @[LZD.scala 39:27]
  assign _T_69 = _T_66 | _T_68; // @[LZD.scala 39:25]
  assign _T_70 = {_T_65,_T_69}; // @[Cat.scala 29:58]
  assign _T_71 = _T_63[0:0]; // @[LZD.scala 44:32]
  assign _T_73 = _T_70[1]; // @[Shift.scala 12:21]
  assign _T_75 = _T_70[0:0]; // @[LZD.scala 55:32]
  assign _T_76 = _T_73 ? _T_75 : _T_71; // @[LZD.scala 55:20]
  assign _T_78 = _T_62[3]; // @[Shift.scala 12:21]
  assign _T_80 = {1'h1,_T_73,_T_76}; // @[Cat.scala 29:58]
  assign _T_81 = _T_62[2:0]; // @[LZD.scala 55:32]
  assign _T_82 = _T_78 ? _T_81 : _T_80; // @[LZD.scala 55:20]
  assign sumLZD = {_T_78,_T_82}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[FMAEnc.scala 37:24]
  assign _T_83 = io_signSumSig[9:0]; // @[FMAEnc.scala 38:41]
  assign _T_84 = shiftValue < 4'ha; // @[Shift.scala 16:24]
  assign _T_86 = shiftValue[3]; // @[Shift.scala 12:21]
  assign _T_87 = _T_83[1:0]; // @[Shift.scala 64:52]
  assign _T_89 = {_T_87,8'h0}; // @[Cat.scala 29:58]
  assign _T_90 = _T_86 ? _T_89 : _T_83; // @[Shift.scala 64:27]
  assign _T_91 = shiftValue[2:0]; // @[Shift.scala 66:70]
  assign _T_92 = _T_91[2]; // @[Shift.scala 12:21]
  assign _T_93 = _T_90[5:0]; // @[Shift.scala 64:52]
  assign _T_95 = {_T_93,4'h0}; // @[Cat.scala 29:58]
  assign _T_96 = _T_92 ? _T_95 : _T_90; // @[Shift.scala 64:27]
  assign _T_97 = _T_91[1:0]; // @[Shift.scala 66:70]
  assign _T_98 = _T_97[1]; // @[Shift.scala 12:21]
  assign _T_99 = _T_96[7:0]; // @[Shift.scala 64:52]
  assign _T_101 = {_T_99,2'h0}; // @[Cat.scala 29:58]
  assign _T_102 = _T_98 ? _T_101 : _T_96; // @[Shift.scala 64:27]
  assign _T_103 = _T_97[0:0]; // @[Shift.scala 66:70]
  assign _T_105 = _T_102[8:0]; // @[Shift.scala 64:52]
  assign _T_106 = {_T_105,1'h0}; // @[Cat.scala 29:58]
  assign _T_107 = _T_103 ? _T_106 : _T_102; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_84 ? _T_107 : 10'h0; // @[Shift.scala 16:10]
  assign _T_109 = $signed(io_greaterScale) + $signed(5'sh2); // @[FMAEnc.scala 41:39]
  assign _T_110 = $signed(_T_109); // @[FMAEnc.scala 41:39]
  assign _T_111 = {1'h1,_T_78,_T_82}; // @[Cat.scala 29:58]
  assign _T_112 = $signed(_T_111); // @[FMAEnc.scala 41:64]
  assign _T_114 = $signed(_T_110) + $signed(_T_112); // @[FMAEnc.scala 41:45]
  assign sumScale = $signed(_T_114); // @[FMAEnc.scala 41:45]
  assign sumFrac = normalFracTmp[9:6]; // @[FMAEnc.scala 42:41]
  assign grsTmp = normalFracTmp[5:0]; // @[FMAEnc.scala 45:41]
  assign _T_115 = grsTmp[5:4]; // @[FMAEnc.scala 48:40]
  assign _T_116 = grsTmp[3:0]; // @[FMAEnc.scala 48:56]
  assign _T_117 = _T_116 != 4'h0; // @[FMAEnc.scala 48:60]
  assign underflow = $signed(sumScale) < $signed(-5'shd); // @[FMAEnc.scala 55:32]
  assign overflow = $signed(sumScale) > $signed(5'shc); // @[FMAEnc.scala 56:32]
  assign _T_118 = io_signSumSig != 12'h0; // @[FMAEnc.scala 65:35]
  assign decF_isZero = ~ _T_118; // @[FMAEnc.scala 65:20]
  assign _T_120 = underflow ? $signed(-5'shd) : $signed(sumScale); // @[Mux.scala 87:16]
  assign decF_scale = overflow ? $signed(5'shc) : $signed(_T_120); // @[Mux.scala 87:16]
  assign _T_122 = decF_scale[0]; // @[convert.scala 46:61]
  assign _T_123 = ~ _T_122; // @[convert.scala 46:52]
  assign _T_125 = io_sumSign ? _T_123 : _T_122; // @[convert.scala 46:42]
  assign _T_126 = decF_scale[4:1]; // @[convert.scala 48:34]
  assign _T_127 = _T_126[3:3]; // @[convert.scala 49:36]
  assign _T_129 = ~ _T_126; // @[convert.scala 50:36]
  assign _T_130 = $signed(_T_129); // @[convert.scala 50:36]
  assign _T_131 = _T_127 ? $signed(_T_130) : $signed(_T_126); // @[convert.scala 50:28]
  assign _T_132 = _T_127 ^ io_sumSign; // @[convert.scala 51:31]
  assign _T_133 = ~ _T_132; // @[convert.scala 52:43]
  assign _T_137 = {_T_133,_T_132,_T_125,sumFrac,_T_115,_T_117}; // @[Cat.scala 29:58]
  assign _T_138 = $unsigned(_T_131); // @[Shift.scala 39:17]
  assign _T_139 = _T_138 < 4'ha; // @[Shift.scala 39:24]
  assign _T_141 = _T_137[9:8]; // @[Shift.scala 90:30]
  assign _T_142 = _T_137[7:0]; // @[Shift.scala 90:48]
  assign _T_143 = _T_142 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{1'd0}, _T_143}; // @[Shift.scala 90:39]
  assign _T_144 = _T_141 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_145 = _T_138[3]; // @[Shift.scala 12:21]
  assign _T_146 = _T_137[9]; // @[Shift.scala 12:21]
  assign _T_148 = _T_146 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_149 = {_T_148,_T_144}; // @[Cat.scala 29:58]
  assign _T_150 = _T_145 ? _T_149 : _T_137; // @[Shift.scala 91:22]
  assign _T_151 = _T_138[2:0]; // @[Shift.scala 92:77]
  assign _T_152 = _T_150[9:4]; // @[Shift.scala 90:30]
  assign _T_153 = _T_150[3:0]; // @[Shift.scala 90:48]
  assign _T_154 = _T_153 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_3 = {{5'd0}, _T_154}; // @[Shift.scala 90:39]
  assign _T_155 = _T_152 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_156 = _T_151[2]; // @[Shift.scala 12:21]
  assign _T_157 = _T_150[9]; // @[Shift.scala 12:21]
  assign _T_159 = _T_157 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_160 = {_T_159,_T_155}; // @[Cat.scala 29:58]
  assign _T_161 = _T_156 ? _T_160 : _T_150; // @[Shift.scala 91:22]
  assign _T_162 = _T_151[1:0]; // @[Shift.scala 92:77]
  assign _T_163 = _T_161[9:2]; // @[Shift.scala 90:30]
  assign _T_164 = _T_161[1:0]; // @[Shift.scala 90:48]
  assign _T_165 = _T_164 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_4 = {{7'd0}, _T_165}; // @[Shift.scala 90:39]
  assign _T_166 = _T_163 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_167 = _T_162[1]; // @[Shift.scala 12:21]
  assign _T_168 = _T_161[9]; // @[Shift.scala 12:21]
  assign _T_170 = _T_168 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_171 = {_T_170,_T_166}; // @[Cat.scala 29:58]
  assign _T_172 = _T_167 ? _T_171 : _T_161; // @[Shift.scala 91:22]
  assign _T_173 = _T_162[0:0]; // @[Shift.scala 92:77]
  assign _T_174 = _T_172[9:1]; // @[Shift.scala 90:30]
  assign _T_175 = _T_172[0:0]; // @[Shift.scala 90:48]
  assign _GEN_5 = {{8'd0}, _T_175}; // @[Shift.scala 90:39]
  assign _T_177 = _T_174 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_179 = _T_172[9]; // @[Shift.scala 12:21]
  assign _T_180 = {_T_179,_T_177}; // @[Cat.scala 29:58]
  assign _T_181 = _T_173 ? _T_180 : _T_172; // @[Shift.scala 91:22]
  assign _T_184 = _T_146 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_185 = _T_139 ? _T_181 : _T_184; // @[Shift.scala 39:10]
  assign _T_186 = _T_185[3]; // @[convert.scala 55:31]
  assign _T_187 = _T_185[2]; // @[convert.scala 56:31]
  assign _T_188 = _T_185[1]; // @[convert.scala 57:31]
  assign _T_189 = _T_185[0]; // @[convert.scala 58:31]
  assign _T_190 = _T_185[9:3]; // @[convert.scala 59:69]
  assign _T_191 = _T_190 != 7'h0; // @[convert.scala 59:81]
  assign _T_192 = ~ _T_191; // @[convert.scala 59:50]
  assign _T_194 = _T_190 == 7'h7f; // @[convert.scala 60:81]
  assign _T_195 = _T_186 | _T_188; // @[convert.scala 61:44]
  assign _T_196 = _T_195 | _T_189; // @[convert.scala 61:52]
  assign _T_197 = _T_187 & _T_196; // @[convert.scala 61:36]
  assign _T_198 = ~ _T_194; // @[convert.scala 62:63]
  assign _T_199 = _T_198 & _T_197; // @[convert.scala 62:103]
  assign _T_200 = _T_192 | _T_199; // @[convert.scala 62:60]
  assign _GEN_6 = {{6'd0}, _T_200}; // @[convert.scala 63:56]
  assign _T_203 = _T_190 + _GEN_6; // @[convert.scala 63:56]
  assign _T_204 = {io_sumSign,_T_203}; // @[Cat.scala 29:58]
  assign io_F = _T_212; // @[FMAEnc.scala 85:15]
  assign io_outValid = _T_208; // @[FMAEnc.scala 84:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_208 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_212 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_208 <= 1'h0;
    end else begin
      _T_208 <= io_inValid_phase2;
    end
    if (io_inValid_phase2) begin
      if (io_outIsNaR_phase2) begin
        _T_212 <= 8'h80;
      end else begin
        if (decF_isZero) begin
          _T_212 <= 8'h0;
        end else begin
          _T_212 <= _T_204;
        end
      end
    end
  end
endmodule
